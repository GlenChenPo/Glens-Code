//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
o3rKLIJrrI4PYEbKsaIvKyZiHTIq+wGchaB6ZtikmgpKloWiZ3vRuv0gSFK4RXM3
JF9YF9KsASqfcUSDTO7pK19Eao33NHC5w692z50KdJWhrGkFwKeqxOU3e44Uowy/
V1RWfvgHtqPLBn7dXhSOxoPKQePa3ClK3X0sEFdfpK7T6xvkaBIPzw==
//pragma protect end_key_block
//pragma protect digest_block
El11LYH0JAigRO+h5YJU/NtKUIo=
//pragma protect end_digest_block
//pragma protect data_block
uo3NApABGaV9pkc/0fDiXrxaMPDEm9KBEM9dJyFTqfD91yf+kKhUC8KN8AuQzIie
WTA8XjXFu7GspKapjK39lDEY0qGKG2SbCxx3fnGNv2iDFq+BDNK6PdNcxO82a3AO
ekuYAlYiCnHGA5DCXRHQvgwICB5Q4xuVBkZZyG0wDHfvWxxc21tET20lIcaW647U
JldMaQzcR3/aCLGuCwMpbgkboQXl5SP6Ws5eBfZ5kiNgOD3tF7K/m2uNDtvJejUW
hHIz2y2TNnW1JcdD7YiTZGuDNzLCwmkjBX36t0g7iRJn5uTQdJz0sQdvj4OdeNs+
FZiy+/NKFKVAXLm42URtTw==
//pragma protect end_data_block
//pragma protect digest_block
bRnr57RpM+762inAhWSyy1gx3m4=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3f9eOiZGg8t2jfoVdFQlxotTSqzdckcXlrNNAuHaVlSJVua1IKvKSy7tLm16O6wx
fweS5ngw1s13KO+EuQlQI6MGY/lJC7T0AfBo7yCemoJeUV/aYiF+fTnwbyfiEIo5
O5PDoCnMcGrEy4oHxommFAup/ArbHYHv2oOw06Ow/gVefEKLEtWTZA==
//pragma protect end_key_block
//pragma protect digest_block
I8eK9LMHvi87g/12QUGj+appd/I=
//pragma protect end_digest_block
//pragma protect data_block
2wiJgoZwO06ctWwmHdoLpmafkZO59o+KiSAWStC/HySZ9u9swyUf7rLvMssuw9uz
sUAH4B77giyQhIIELb+SPhHB4ynL/AnR9zZVWf0noisr8BS9KUU5iey1+OnOOPrX
GdUV6RQE5TGny0kn+CnHvolTVuU1slL667sktfW4Qm53uHSm1mgNIUm7OKDbjMlU
pZvc5NwTvALKz62+YM64F4mbJCA4DwTbPtiQRqHZpe+TD+VkIFQbB/Q0kQfoLlgi
0xKrJxTUSyieT/NymGiFnZsIB5KTzDRnjNGeWc957xBKWMpwH6omRofk79BJixw5
iRXxRmjgWW6+Oz44xnPBdQ==
//pragma protect end_data_block
//pragma protect digest_block
9lgR/5/DUKt8rTezxIgoHOpC8HM=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7JesjcHCMOwVASwsdEpSuOpN7nSfGuT9pdqkalbPf/qV3uVMtQGJvBUN2JOqLXoo
jG//z5MkSIMtosb2mjxf+507/14/tJchWfre0It+X6//YzYBaUJXy4fyaAjCn7dF
byTDrjFTsvT0mV77zbRZT9tRzmEAUgtioYeYajKPpJHDn5X93wA2Kw==
//pragma protect end_key_block
//pragma protect digest_block
+ywx9Q7XgbI7FZGYJEibKI2rpSY=
//pragma protect end_digest_block
//pragma protect data_block
W181g6/UhToSoEzX8xEa5yoCG5brtO8ex4gMNnciv5tQqz5QDw7xzRlU4IYi1pYB
5E+0kAFM539kpuCdb9HcTHAfIVUWHCP9vBgXIt8FISHOMBxcpBIvHyM2ofJaM5Cn
hVVcaQbuaB0PNtlgRxj04YDNtDhlZ6ytBgsSy/vKV1umg5ErKMGWuBfhtsHW7ID9
6sYiTo8ra6BiOq6SqWCE/8vy1xbCdkRj1BPs9bj781ZK8i3PuL5LzI3JKOwvlFLP
nO+9FBItU1qoy+n1twtZ/YmUCmaN7XbN2vbJtJCbsP0gymPc7hg05aFMcjKPTii4
//PrGzvi39JwpqDy/9ywztsl6G/VA6OSWzZXGb/mVqf3UUFDA8yi/NLoAxNojmWX
xsKQ5Fa0IDIZoQViKe7zbc2CrUqi6g39rtR1m/gRpxLlR4alq5Vm8nsuVqPZJpOo
3iOqSGufutvSW5x6LJOVRDhX4FMzROpT9nrK3q6JLNCjh50zTaVuRjecpzZ9gVIC
HTC/EhNIdd8zAtET3bPPFXonM1zDD+rqRsu8TuXfW0v0T/8AH4fOiWrpDKz9u3Qb
TeZQoADLCPUjNYdroEK0yzmP4LcMGfvsyHfhrsXa+wVu/gqTVYhtM8u3v+RFihoZ
qChJljs4wQcryhlw+UDwTnjMJ8wY7glrSuODD55aZet+St4kNvXkDjUfdO2yAxCb
iMnJdZ1sTI3pANC1m05RNaaxVhcdsSeyFLYGpDCOwkq8AVlfMrwzOBHu9xPF8cjP
YvRXr5dXiiXDIEzcTxMSd+OSqfKuaGc52wqEnCobHc7h43p6SjV3tc0Y33v4ZbNu
fiB2zGSMgHxEIkziNSZ85yQ+HDeXbsXcj0dqQzYvuchLuC2IcoN0/UHnD+HfjrN1
/g5TtNKC+ztPw14VOeK80iudgIpB4SGvy1Kh2RCss03iRb9TUs7O1378H032G5bA
J021xDhOGYIx8ScxyqWoTHD4f52W/HKnsuqCAIXwkBhzmT9I2gMQ2R2lur5ZQeoE
aD1ge9/Eup/si4dx+XinGK6gIMkOnTK9cLBkLbzn/snfCkQNRBfJDBdljPRYLu0l
xfcKDyOPzDhWtk4v+xS41qLhgSS6W5Dan9fEqeV6Ed7t73VL+ecwC8U5I2GcBTS2
ZT62B/fJUXfUy2u+zRtjtzhkpLx3s5EQeDLLj66Vj0kcg1dMQag+CJ2fEPkLWnvr
Vm+wb61jnzgC8bTX489Y3DZHEvyE4+R/UEYHwVY2bFuRX0AgWeZVDuPhGhoeTpzx
diedBkdszLfA1PkKFj7tOaEONNDSMj7buuoumdiHpHXvjDz6UWEgCAP3gFpqnYho
0iHCkQdWPC3uCYmrFDGVSVR6HVIIlJupcbsUrzkIBLQcGzrTRI7vz/IaGapOW/zg
zdqEwquhBMb/AmMkDaxU2MjMjfwhI8IGgkaW4n+KSmCYm1ryAUlL8JLSD3QwCFTr
IR7YED53ujbPzuZEOlkKeGTv8TkfS13SQC37JFOGEiQcbcdpnoCH9jIuraIYlrrs
U1fPmaWftuBRSP3XNxAyFgqD7nqjtE8y7tvWOY6jgjd/MWFPBk4RRnohIFvbsqoI
pQ1FfLY9iUoHAla6pW+R10xQEMqnHHP3shYus02t6TidwVe8IoLtRuNpa9Dxx8Kp
UJ3hwZ9f9L58MrKKLg9TF2WvjAFoa32lUmVbGoHC95aWitcmmRTTXrn8wRcAnj4h
juBkWWliOiarKQ8yEXAOlb7tvdNvyMpuFaiHV3PEjfITurQzpJImLg1nk6cLAD4l
uD1mUYuii1KOvJqc6pj3c+sQtc8W7ClulNJ6k3t8hWx2NAskvAwr/UrT1LMjkave
jjADL2qn66ceif1Ja2PuRAUNLymFDkfVTaIHtE6nOyAXnWZyeso+gbK1Hbr6tRIT
81WwrcHFDBQkVKKpuCz7QMu5ovs3nFDwyba9bX1xM+KWIM2aS+7oWmpbQwFoNfUf
eYoEmGGBWOSVooMK5FXkLyb/TRWSke6LGhAQwhfXliR5huZfct3XzSVpxS0l8kqR
kW0SUJU1SFhCfNbjeGDI4M9uHJsoT0SMkihrU01towlK3hCmVzITt3cNkvzmIair
2CVyuRZqWkzDiLLX7hCH9r+SWc49Hvb2VL3Ba6TLZzgtAxTXJqVRXASAXEibEmnf
4dnNAzmWtfC3Od3tsDFCl5W/UHvEP9FNPZTEVcOe/u1Y79zDqv4zwfk+ARQCNjua
qwF94PAfjlWPLrhChuy1Y8yY7LpCvz5Yhzu4F9O+elnpmPq2qXe7MhvuEfUhCgWB
eJdS7sgnVs9Pr6FBKhP/bEoliA1Kw0//661pGzrKRJUIBr3sSF/RvNtD5QCIEpn6
mRIyKNB/PpqntrVhfopBV3VfaqJI+M/Q5UkfHNoNoL/J/KGIFuoIliQAZZY2VGEL
L6fb/skHvAB1JHVc5J1xsdYkdTXAqZjoYO1+Kt4RYzBug5I1HxO4zqr9NZCFD51r
l1WsL3I1u69PuOc+ALu9+6nGoUos0USbGpi8wLM+gFey1uSWIDkmlgl5IuzaTvlr
iD+z+LgVxQHY2YbrEVOQAwpe9z7mz5rngqZpVNdMHa4XSFJIh+Oanxo2p0otXGhN
BTM83sXp2cGHidYAeBK+be5D7mwJHcPiCYE0dNyOmKfoj0TdN+ic0i1gRK7D/YAV
ONpfBwzK7PUoAgSaDMk5NB70rd/Ec9cGLg6cmVIAyDum6jqA/1RDYbIArovNelMR
5pSN2C4TEfE5StZrJ6Gst6+RvqU5Y+tKLcxz8AvJ9SLC0w8Hc3hCZ6JfBxR5zkhX
wn/GBG90gqsnVcZVvz1AZ0TdhJyQlOJHuokO23GXoqY5cr3t70MVDPEf+OEKu1TQ
uOfpbyI1v6PB5gR3ppPFItoI8zalxfJWDQ/sdROmwuiVMDms/pLYuTMCnEG80mKj
2DvqKBoBSQTsThte815yBsJnRzTdi/IRALYLMcCKKsF+7+4kkIKvjjqoHzAD8XXp
ObZLPvZT1gQN+FrH1ju6JfNr9zbyfYFKAURCGwFbiFNRPBNvW0sp2oXOQojHSk0p
UbHh7fUEjehVaudpeaKaCRLFlMoAZJJHOHtDdLuqtf1uI6rgLIBFIsq5Dq4eYyz9
gsAbQZTPgOCI7rpDUNFi9XDYsrS8U9/o7fcc9In82mIA/SI/zlM65hHFLBjfGW84
06/EKtuGTmQxTM7C1hm0+WPj2jVaCRSTMaHKfv7K3BQAUrbJ33Y7iIg0uXhgsuDT
Qpr4Ut2FxKyILyXNCinEB3NDSC8BhDTO0UOxdjd6JdWmdpuGoB8ynlAefV0qqUBa
100sfE0Kn+Pos3yxdHPS/+qd2xmLzWvAPOjBu/Wnuu9M7uafbYSOQIPZw1qPNfih
hr5NEGxbhD0Tw452s52bUauoAVoQtq495Q+LzAeCyTft8mAQD1M1V3VVD4sQ5Cpb
lhEC0cnWyxWL9l6+WL+1owlv0AgV9J0nSWLUfH8MApINxLNC7ZXtUeCinV0dImVp
3LlqQK8jMJM76hl+Mazz5mnj+VqSLQbmJc7J+AIGXROsXZBQbDopfq3V1CUzy3xl
DfLC40R6qVBNZ7BjSdrG6pnscFgrgYowQH08m2XSg95TP26s45r0gD2i+/Wqkne8
zH7Uu7f6U27Zj6iNxPPCiG3LyiXd+R3ysGZgKqaSzLZzdGWwuCUWG2Iiv36uY04v
97nNKotyr0GmgSslReYVpTNhWxim6M7ZI89PG2KiURqqKqAMbiiP0CQ+ajxm+to6
rukb2ya5yDkriLCmHHwLgzmxOQuQ5eX8xSR5AUS4cAyXJ82U+my6HZWzn9ykWjaX
Fw3tBx9+ThfEyUG+mdICLSPi2jQlxgxkFcZHWS7NYGVY8u2g3xmlWzRQFUSENGiQ
+9atqmkdf4ORe+kouhcZDg2cKYp2qcxIMk+/wq/k+f07kYC3CbEZ2m0BsnXN969x
roJwqMrecAjLHX2XFESs33qYN55IH/iyCsJTDKSO8pYdzYkJUuqlw12fepsyB0WK
Qpc/pwsultt3tBkc1h7jo6w/eMIsilES7FrL4loLEJVHhJY8gael6M2GU/uqxVD+
iJGcBZgHRrPTk96TWfdLEbVs+bChkpOreBDglJBdPzK4tl6ou+Zo7SvOz+HBStbc
6la/dDReAPGkE2l/ATfNt1cfXxWrWoAAiupuvMv6CbJhfFbmKgryAGhSejoN/KxK
whuLZEYpGAE5gWW9QARMZa6uaxdg8QuLWGdHg9GrYStx/jAK0CMgOTCFvMaJ7a2W
RHjxXkvDEEGtCLjJWee/BwKdBOvuB3o5Cch0KaiMApax9A83P0EoOBTI1GbPXhFH
3szX5qszmcSiX+RSfLFYTY41WbNCD3UAaZokl02cxZN6U70IgayjTQ6ZmPSmH3PL
xNaET16crychfvX2n+VChABaarVgTo7bef7X5RsH8IDVDWa1MUfPcrCllwKm77oq
r6D3xQzxBeUc1YahoXDi3fzdd4x2ehkD0QkpanvroRPNLIK5toBgGwWh674Tah8o
WBX+fmwJ1/sZpciDp81V+zTZfNaZTm7F6gQsMDJRrJcKc/XeU2XE/v6RzOs+areI
qkHCVWR92gpWVQU/yenghKIvLhMjgj/hLPlGFYbJd1cNj4IMd5sy+ti48tflow3f
IHdhYUVwOfw52gIEm+oFxtUeHf/R/8LSvPyZ0WD9wBznsE2SBJHjU9QUNT/nDvt/
g/k4aoPxBdZKNbjQLtg63tU8hQQHb8NTsgzelp5tH1wyvnhnDBrnAo/O9kXejG3G
9k5ITez4l1NGT5BC+VEkpKXLke0RH9F8w8kbXhJKVTKTh/jc0dnsb6SfuWf6oEkY
LECNg7olynvlioJODjankxUJ8BhxSX/uHxyIACy2VPKuWDJH1ZhwMIJaAUxU8eCY
A/h/5owT207xPkEwrsY3Y1vm0JW+++iasl85boFAk3sBGtVGLFeYHWeCHWrjXPgh
PLq84idWeDxHqw3ycpHOYezu0rsJEEaKubsEKc9xU1+azvOF3+634yJ2se1nPYFG
OEl5p8btui0p1eAPUoxihZGGOEIn2ugDtm+ZObJtm+DqiyDkxllWubYL6W/XoXiP
FtLSG89LQQKXZYpQ95cZTTjw2mPWUODJZj2tcBunAQ+9O1jkb+UzgF+/zP0ZBSbL
+i0Up4Lftj5sMrsuPbSOALrdcWYHQ+RwLv1blvfj5M0AEiGc1m18RBDoQTPexEzm
lLQ50n/dOt2zV1d/k2/4mn2eDhDPfZFOIhA+lE7UqfwHDjeSaSNeb9BvfqSC1h//
WccHWutvAgQYlN/uaGqBu+MhcYYWPqfUPn0mDM46ho24LvtnK8c2RL6F1d7qI1Au
9yyrbbDkUbt+sMdbMTovvERykzsR63zoS90Pa4BJUJYY4lhQseKz1bQ5RkhzeySs
Lw5D9fU1T/M65/BCttOvz6yPB83dJ4lxMM4/3w1yU8G81KzXaqpZYuCmqFSP7k5E
ub+uxZx1VlNVSZmnqQ4RRtpHOPcx0TFwEqmKBODUSzArZDwwIVC0oq/KdcQC7178
j46wstPw5TwKTVhrulevI9a+5CUKTDrNiCYLNmnqN81Rsf3Dr8UiesfRXlGZkBWh
OAuWGusRtVLQaZnc4WMNEI7bmwIJztFhNcLn8hpLpZyiudMphrfzdZHRRkk/bCif
VUWq6lPDtJvi6KWx9XB2QuVQuDWzomlniUJZ9/EqVfY4lgo3HBskkhi1RbMJJkBw
Xb+8CyGIw7GkJw4RZChh1ErKaMI/gO5ixiyygjvX5alo+jgyinJRzVNWfSNjLOQW
8hvwROPhzBXqKlI8nPw99hu+0AagUM0xfSMseY35EnL2J4Z6+jaYtb91r4T9rQf4
W2E7zHq2ukTfaRjpNO77NiXpN1abinAk6bIerEvS5KKjaRw4YqJXAG9H6zNG+dcG
tniQMBRwULadwAyJrcwbxLYX+iKV7QM+PC3EfL/Uq2w/TZOrtEYPuUSIw6FlES6y
GCI5xJzJBMAUCx2fQBTJ4XGd0G0fMVPi1lAf31zP5seieVUKO/WU6B3/V9Oy6IUP
tfXAoiA4hhHwIOZeePkgk0gJRoGRQ4RJ8Ixz7/JDfWdvouySDmIPY3YDbD4G4Au5
UTH5b8nNbpqUx0kWdYHr5IpsGSkFyctKyM2lAlQQQp5caDYGhASzKEHzGpFCvT00
Z/ASJHictd7ENJFLSO7SsCqX738vCHML1ok74JkCcAGTU6v+mbxR7MOYNyPVILQK
qO/rmE04ToFaa4RLRn7zJkwuXZelltQkOrVif4g/0wkaodBlRTKlAUAegMm3T0ID
/An4qSSR/Jdp4ddsqe4i9VFi075htSGGJOBla6r9gi9EH3iJeRg+Oo2CY0v073kT
JA1RLIZss9N1edJcDUukqgP4Mz5Tj9Q/SBXp97C3KdXXaJWyJxK3t4nbc9noeRPL
p4ZrZsItB4rhJgbtsevQMdzp5LKMuy4zf9tLSk/4Nwejy/Zj/D0ZvLwx554ey3rc
6UajCLEzarVpk19AwfrY6UHgfV+Fxnl0bjNzxK72MyOIxwKL+uG5xg1GJDdgyy41
EJnNiGJqWjrb4KNP2F7lzmMqfC2J3fCkYoHBEJxcyzpzl/1SXC6aBraEoLIL2M9H
J46e1OkcDLlTHf+Y8enpQaIfVbyjc24j5UVfdDvu6w7hN26g5Zx1czsan424s6nF
qd87bqxChTKey4ZZNdY0dmo85lXDtrIFIEROTRN7YBrogEEmdctm4W2lQAWh+gce
cab+YV72WKPp+pkRrbzOjWSpb1CatXNa/Rcw4ePfcDyF2FG+a7HMe3WkOWGi9YLJ
eyEOVqXND4LiKkqZfCEtqrcIuYxuIhzYuDQV3bb+ohWbiHVyq6ialUcJ5Xd5i9cE
Amu8r/DZA8pm8KBNj3v6xrZGW5+90RF7fp30Q6Gnmdj+50GHQ8qMUTco87CpcNOz
sbSDS2GQyGfBek1BeSY+q+DNQo+VABZH7S/t2Mpa86Yr1oBfB36uSpL2Zoq/0y7R
JkJq1qAaGhlS2D6rK5Xg84rm8JOEQHQPHemSw3b/zhP+OT+l+ccO8UtLkmGp/31q
iriUa8L69+vMVlsA7QcRVFj79FApwEc/r/+CEPArpyYHKn0ujXj/bTPxkRFgCH3J
USr0cfY+NbuS/c1skEzUYw5Gi0qay5mzZjJa1S/iQL1CIWAGfqJMhzK+0nLwoJdb
vq2ISoGSOac2GQfoba7rB7ioRow9ghvGjyzCiLvUkdFedG0kOKlxcqOO+G0H4I/a
FIZ4dDx8fMSJPiFc2/N4R7egmpkOYq7AG5bniCCOFEe8KOiDdeaGfBO/ThvAeLOz
JYPPBETG3An1gK0w+d1fVoGaGPWGMOfAOceXrQNLg7uoex/wdoZv+8COSHsGDOma
6+IJ29bg/k1xQMTy7IYyoY9ok6Yp0m58d0RV0r7FFQdUSZmeoU2MHIWlO2LNSG9p
o+LbwJcZ6H1zRvrV+IsIZl2Q/Qu2UbeE7zP6mfbOFMqptqMcCIiEXWWgeepAjY6O
iVPZOav2+U7Ff83mB3/hr6KMqNZoES2V9fqHVdTtQVHiqPJNWaHQoiNoVkBY+hhz
LQFPDTcMPcNMdvQU8Rm9mnHQZKqzvW3NG47reka14egM0xKDJ431HATfs4ja5IlE
eIQ2zp/h9AOLBvKxbckpqKoq+8pwxAO1kFSYFsq9bzWcYHp1Oajp30YnQgznf/lA
1ZLLcdj3qXn9IUT40kIIDwFc4fm6IvzPvBmDiQoloqmKPZ8ckzoG9wrO7S+nOI67
zwdf89kVbJviVGSkwq3KDGV9IRQASWUVrY9WZRAtlF8Ij6WYWG5unBPlZeo9bIwH
Rb7iNG3wHkNSXPsWHLkiQ8I7pXGyCow9K8J0iQWXMHxIRv2LHP632qKrBUCa5u3C
yB/13GqqHAQIHyHoDXN/VdFrBoxLGZ9auPInAVy14K3Jy5qi4M97WrqKJf8AtRBi
PdrTXCmOPmttS0lqRtl2Hgzacih7OV4KKTyHe05huyidc+TN0/cn2bKWUkIPtGRY
V/W3fTLLvWpuxx2cdLMsS5h1/hCgXYfpDRACUU9bRTIQlUwHAV1d+R1eziqRfrHG
rf5ZvPjaBj7bMvwve0Ex2G+0XzXAt4GFL5g7HQ5NMIezPmYuZMh7iKdBKeLT1azP
icTtNHtEPkT9aIULmxj69Q0iT7Zn403AC/rszemwvla/DBf3C6J37qLmJppvG9Nr
Ao7NDZBKxe/g8wMal9kfnfemWZeBvLgus97Ft6HiBVGLh+S96r+Y3wh3Z6WVODej
dWe7qkaCW5/uKd+S1xa2kTQpCkuQMoSTJvO1Le2ZWb6ynHoPebH2MNrGEFbvZSZd
H3j5oHsUOhQ0pTmUL8WqkCeKt4vTWEsgxcoAKx5ZI4v1DS4+NFqtUa7xg804Zgkw
g4kRUQKIBV/SwO5nyNiIZv3aby+AzdW7JKbuSXUun+EZaDZzMyoVyie2KV7uWubR
z/7a7Aave0L2b+tSDyp+7PgY7SEOomcrr9e9cTd6RrOIRnhEW4EBQEFYeMcjNkb3
JFUqfh95b3FWwksYRrNsB/oSiI/eNVv5pCGZHyzhjs587pLRtW7ghtqjJtNW5AU/
yYbWju8dLkFGZotqMYiOezoAmTzLD23Wv0DOh4gixWylevibB/9r/oTtkDM/+dms
ARb7Tpuluy7KVaDj8pyqlSKAX8f+7VvEdn6gyG0YHDpnLu5j5JEObz0AKw0r3R1m
06NtMPwZ5e8J4pk5D/3VmLTV6AZieJqAKFfSsfB/ladl1sLfnazs7c41ut81zdG7
zhuIv+ltceHlbEUlUHp9fhHpML6nVhLlsm+oikcZ9yEDzmwP2Hh6tZbqTRNplJXK
PahmV8U8HqBnUAZuopnrKkDe6dn7UnL1X7G8FDwnZJ/2xzAOV/xO71Rljh16Yx+b
p2cr1Q7rCiOcwQRIAMFJljHCLgNAi1dcZQkv+6shc6w7+7z7BU1kcl+87AdH/yhH
ljFdkTZqzBU9RoC//4KO8CidqKcQo2oBLNx+rLMtQB1dYHWzYIm6vqeHsetek4v9
VnHZVpZkFIaxvtmeSvrfcuODRZTeZPfRTG0asfuYIPbswYnu7/AhyEt24JJJYi1l
t8OefOEsLvL2eORVuUyFLI9n7Ip4rEmRYATXvJkDnWsCrOr+V0oK5h7l2mpqEeG1
vlVjEOUG8efcE3EKcspLV3nzJD7EnOmuLQuy3bM3WhINg6r+5Y/8azPEK6ajCjRH
s4wwGKdRJk38jqvA5w4ARgm6Q57PFQeSzih5VAajisDy3FwUlsJbkF2+xF3F/MVa
5W6hkOMXXNc1ol5Afd8KLxQtKbBLZ2mVKrfWPvfRbjAn+k1J7EW58llPS9Z960t6
pzdomjNMyeKysRK2yH5yMcv1ngdUVWt1jD6r6bs8Uq2c5+s08SQxEYm2hNLK4/r3
XK9e4Wu4FHMHc7Fqb0aZXuh2KPt0wZDcO9wrMSZ/q5hZ6qp/H3Ye9Ist99PXnMpx
4mYKgXbamfu9vF6s4/Aqb0khw4Yb+ZtQbY/zJc3Ixouj3VRVmrkUZ5/s70ffy55m
lPX3ZSXKq27towX4DCLjqVZLkX9LamL3abEEk8GVorLJM+Q8nVEIX1NyHe7XTlJW
Qv0R1AJaIWuPA5mmYQwB+KPopyWkA54BYgqeidK+bH6n4n+RTMwCyTPSAOH52yeK
ExrlFTWzo1zy9gOjOuwwF9oNAkOAKkTHLGRuiaoqtTAS1WWGD3jdOZPLHT0Q+2dt
C/HiqV964OTcQH98EirQfRfVQb+/99cHSENdnXvqO9bzqAq3t7u2oMMpVH/BfJbu
4b6IRJ3pnGm6N6A7nOqYd0bLco+aWsKkYO6lVPfhTc5h52R9eigwp6qgGUaApaMs
IRFtUTI04r/ULGyv4BFhRkF3aU1Pp5iFFP8X3tNou+NPALWvocUYsO7YvP2h06+Q
ohZbPpfSbCDG9T+q8xTfo/Lo8O7o7M+PuasTxXiqVg96u6mdygF5nla9QlN3/XuH
QUS2FLlB6X6VhKB90IOl8Q5isSjgQxMtMCuq6t84NBckCQCLc7A0v1iDzNnt44gj
d/mo4dsHMQByHpXRxHbj1/X/QPl1Lx4pWC+c1kzcosbcoA+QdcqHuBf22guIrB/A
eHwRp0OudcP3yViRAmqra3atwY3MSbWGR1eLY44tuuhMq3b+467xS/5cYm2DECi1
04HzIVVAC9g4kiv58sjO54+kxMr40D9YuC2l5M6Fsq+DHIEfE1w9HN8GrRNqXLz6
n4JC3aWcqwZZjhnkstWgfeqL5HrPI0/lJVxB9YbDgdZnYEB3b0LS/fGpNphdvg4q
oIzW+1O1eS94Btt32sU+gr5Msu/iawr4phMdZqz3d9J+cL4TM+lrzvg8lmBBmNO3
3C1zq2kmmih1/B2a3f1gWzIf8g3ZfaavapmaiShTYfp1axPb/3QtUzEa2TRieJrG
78vglE1thgmAA0YtAhoAU+st7VM01vXBQPrgqSynvAZB1CGLbYA+2/wKOpmA/yVr
1Wluzvm2Xb+LvA3jorkG85FztvCpBHWgyAGcmAzvG9YEi9i3Te86y6EeUdFjlZ2Z
KPhbLaFeWXPbmWlB2voADezNrDuV47qGkSkdaNg67h9xb67OtfK9waZADa16sLAb
JoJ50x455qn4ysKJTZVkE7DoYudB1D/hGZjpDspzuScRXHIzm3WLypD/jYB0FOjj
fISmRU6lyqWy4AKKq5AHPRHrb7JLopL8VatJJT7MJ389nSx6dt+v0s5BBBBoVoO8
7jSLyPtPlxSwgA/Ox6gAbS7FKFro69OnzylagSmL904hbTzAja0zegQONcTvvx2K
ByXwlo9M4hQ6IIat361qdxvvKeYePc02ZqdZYm6pYYCj+640FwD2u/vTrTcwKpVo
Kj1EnTRcRjnTA5FD0rVc3unRhGyVGfY9xpKQBL+PO1Py5qa/zcG5AntKZ4QiX9RW
3IHACVSbuJF8qIqmEC3rIQMB8tIWB3NpBZXSnISWJWWl/S6EOQMGnHBHAWD0+big
f/CqosNUWVGxo34fyhFnpGMCngQQiGUshSM4JmrFpJQx4qSnPG/k17WrwkzJ4pPt
Bq5xjtwoTkAAUFqT4pFChmrM80G+gaPAxLlEyxrq5I20O1PsnAi5onJBhGHGOgnk
dj8+lr962aruSK6bMBnAz5qrMnH2Dga7J0hF3t36pHSWVQQWxpbUfMntZx1mTckL
JJTcz+blTRDRxXLfxNZjF3THnKSfRrDMlARtA5Eyd/UPdVBEM9ZuNqz4wwVe2Yxd
Saq8z+ivydDdiq0GQrMzqlvzA/pXN2rAqoqRE2YcRuskfWwo1pt/FvsgLpSAgkfn
D6s9qW032Px3KOTFQifP7rYY7m9tFmYbIa1CppEns4qao8ePeXF1zuWxPN06/5F5
4vhQKhZxaa4J8fyWfuyARQ9cV797zonETMo7B326wLQwU0u5X2/GMw34AA7pnjsv
MTBlAMBSilG2nWdlB7f7HTiKb+IxnUUIx38fMw4FG+br2hZ0TdlHLwUbn6odhTcE
KarcWcH80OWfYBLE7cqvlpvEbqd3qzdzmN2isjOp2ddHKt4BPTFyYo34Wflyc/U0
sf5eX5F39iAwHsPgJG6aGY+sjJygfHTyprIemeHtLIc3pkwhlQkVDJUCiNKX7JfX
fUPoU2jC4+VhqNKzKYPGfW34s2I09yrYVMwmZ3GlIl6ErI/fd2v7aQuahSoAfPXq
cQsUd7xF8USMrbN/KEkvtUUuOXo17j4dy0BJctqz/LTG/h/JPctNxZhdkSh2wD5X
5ig9gmqcRL4JrnjOTPvS0I/kD+POfi3zRmuQlBmaISsHs9wnwFUW0M6SunfjLnnt
93eVOciG39MtEkVejGbMWmjafu4hhqYlqlcmUtE897X3ebcDFWhuBn5I22PaslwW
NN9mpNFom3/lrcpJt6ap9n+P/1LrCpDU1+y4o/x3HjaTFVLhIiv9emfM9KntGf15
SAYF/ddXYjNQ5DGJxVJwYK515Crsbc11NEHgIHIVccGcTGvemaHxl1s5TIZRiPmc
NABy82bUGNaJwcmz6u8hzCyzDds0N4pJ2cy2xQa1r+ZgdbhKw63uuLBku6HdUQIj
Ojc5HgxCfmJi9Zcra8j2vnmG9p31/psF8LRtNmK1JUeWoXI23PRf1J0FJ6r/rjVV
anRGUKdW2wzStrTbRfvGwSVBkMNN4Wu3RkcezF9/d2OlrhxjaEEXAKr9aTKVlw68
cS808Ofl9NFAeTa8ajwk5+D915k9Qct7wBQc65OlgKZsXysvUPuIBSR4GuPPj8f2
CJN8JuVc0Ya4wqCu7xoYbhVH+B1wsDuOr9YcC1a9KhvBLjsrNjUBQJQ+3zTg9p5a
1aR6Hj+UGtYfWsWdeJ9o3f7pHVwNKX3uAA/LsvBoJY7lPP4PVI6WRkTC+A/4QO+U
YBNfIlpRe1SHuo0HDEOCgvERpUTMyjOtEMWO1YZ2YcnpLFcFrNqmFuYwVi3ZxXds
lObOYL6D6R49h8Acfo1xUPcsEOKzxxKVgCuGWrFqgI/6kJBQSrfNsu3j7nieonUz
8cSfcWq2P8YPBdoQxZ+DdZdp1idcrIdmXeHpH024FZDXl1gumE/aIAMcu0oKW+J/
8V4jPlm/pofYoS0o9p05RdxKti4+j1YTjXLVGXAST5a46IiKSinxeRSBXNbbrtx1
PEqt4JT+FKp5xMMHMGkaYGc4jIEDgK7AVKhOM7o2H492eRmd/PN3egxF5tUkzBaM
VAwy0arljAe+Je373nVXv2vFVKzr6Am1zIs6IRfOw/J2C40LAP39pR6rCc2RNJ6w
dCZnsnbePP5dzB6SIt5dBcKswfAnOeuS0qPRzZxQZtcRtiN9yORfpKcjDJyb3UUd
X98pIpeCURABomfJ9kCHF91cIlMePVAWEos6piA/N/Yfiz8LWWffz+mZMn9K/etm
wYDyMiYSHyleY0gouc73HtiDAzShiSfmCzZVNOFJ/W3oQLSNA+uFq/0Fk5hkt5Aw
DT1OWckA7o1+pr/9UcZ19Xzacf3o1LrlgYfph7sfKjvf6jPmWE1sshsgz1orlV4Y
/tB7BhRNWJKfskKWYktgoFDZqcau5MkWKIp7ttTtah3dwBNB1bamXvHbWfqjYNCj
byBecZ2hYmaNUYrEcZhVusYBfzJ67N4UScqis4DdtHUijk4PBZtbhMUIcsAftfwc
3TaPk8Z5hs53GLhp8Hf0HR63K6D3bYgFi2hbRPNoseIukYq21qPb77ki6wmMOLqP
SuKGFeH2yd5pKsKHogV/pxpqnQ762swnmXwYi7O6ZCv0/7Q2B5XMUSC7q5HhacTs
txhz4SfgUF5ircmVB/DA0F+7FPtQ8EyFi0SQT4XX+Lf5ud5/kJVaUiaGQPwNmkLF
IBs2Fer67w4upXijhUokVCQKvqn+drJeV6PZQmLIf7+CIdf3gcyGjZ7/DV1Ew83t
O2e/RHomNWAH0UFkhKs+cU0OAupvZl+QC5v7/QJjtJzvePlDvRcfCTkhh8j83AuG
WBvH9G3GsoufeYnapieFjQj3UX61+l8EiCm4LKdny0rpJZON/TUv290rm6Y5paI0
7Ma+0uD7lM2OxxTu7jag8M/82sGfI0adXfSa3FW+88u8gXv+4kdPgE63BTaJJRQN
w0Ni2eiRBXMMV96Hnh0tbFpFBae7g6teNDi5yuMicbjnqCFehzfofHNTrQefXEqs
Gzl3LqOvxOj0Qm5BJF2b8dq5bE3DMRt3NoLosyOkWH6jih4dGonFpwlyv0i5uFaF
pKoCxNAcbkVWi39roNTY2CsMauHPNUXE5U1f9ISzB43iweaMr8+UXeyEYKDNDkwf
FI9KqwF367bg6Osm2RnJUpKtGR+z5lqIEpCIjcYA+BV4leHaowS1rzvN8X2KR0BB
mXdjTc6+gLZkRVzBpLyLLHopTSdeTzhTfuxi3b4XzKRmfDMWnrFJU6saiUY50DIr
ipfC/O2vqPJLI5WKoChoK4bUNx2yylB4aW6Tyevxd1NPoG8FZFmEoXbPHkK2wETx
pTsTvTNtpz/n0kNj04h6yU6kXLBGLuEHdz7H5dgvQggcJ9klXsoVw0hGSvgznQwf
3n0S1GeMjMUYeB/9/HDb4EWG6UIFVlIlLZmBDeBkwLR1fwdRIDXdFC2KbLzlEq1P
lGefhXBqU5uzhNykH5BXE4KG7WtyCpst7gi5AIQJiIsD8ioQtFy3q/Oh9B5+AUG8
GU4X2Kq/wGFvBp7pG3SybJtob3b6u2oWYX8Crx36SDdyyFBGIl5wPGa/wNfF+Eq+
YJHN+pxStzf+x02VF1rMyzf57mpoargqKKkP+mqq2HMv1/1edcZ1kzyRfa/veUx5
Z6bp8tijiBmduHViVsHJuYOP3x15O+6CGyZAkhwhLFz9s2ZFsxN1Pt6ZDFD6hqtR
C91WpDyE/pMYSGXEUyXyZ4Yh4Dup4Kh4h0iCxj7N1+zNljMUeb/FB63MZjJob6a9
H++PAc9vap889Wif3t/bEOQ9y5JMGeJ5qXVJEaDbwT+XakFfzcbjyCGizDSI4Spy
ZdpdbUb0W/PkQ4GBdm775RHN/S3A8hBhfNyqpaBD4emPjmis8FO9Zpypv36a79uq
ngzhhgv8sFg29VFGYZ8g+dwFfQxbtTnZ8CrrxTHv97DRRXYNfxtyujrkthYQiWcd
26PUzHfs7hE+JvxZghWuA1nJH+P3zS56Z0yn1Ak26vOGWNpCojhxEVji8L6/BAA0
sATEgve4ARqhoPDxwmsbIC6lK1xe/dkeniXGA+kiqoa+F1hiaY5m5eUb1UMgcR9R
AB116RIBXMqdjbkvD2xM0KzSJdAZSg4UhyRQeGtyF6/y6+WtoRdDD3UPjwdrB9AQ
5WaU/JvxrIHr7gNmDTGrmsBh0wavKgbiTuZU3vQXmemBRPFWKiMYaN/vPscFtuAv
7g8kM4x8ZE/3i6EmzeBtNJOSxOgxzTcTFvk/jaNX4Joutjjqz+It7bl/mJfhQCiC
+oksZ34/fgVBoiuvY8VL+eY/Zx3A4GhBL2EocQn+Gc/d7mXZXy3IbvHDVKXgkt+u
gKiL0hIQM1/SwVMddogt6sfB6qZYb1MIQ/vehH/exu/jNTD7PuEXUQlaWy2OBxZF
NpGxjy59u4t4KT7wFyfWy7iMXQfw7JJ5AH0/mRY0XGeq9IZrX2BgLjmu6z64RqXT
a2D/byVd7DmZGH/t5iHzpAHCS8fqMIybvqMOIwwAGPKE+Dbb9IGL61g12umK20Ot
QHH/B38qeIxKUcG5thAf4STRJ5pFLyV/meaeufen0zliZwyggLkDTZ7cN/5JEVOf
CmPvlWpnvdlpTz5SP3ScTV21gx9g0DcuAmHP2js7FM7wx30C9c4VNyKEFQ5AUzFV
eV1NhAty6Zoiq6IeDyEEZqsv4OYDDBVaAbWYPV/okjw2aLO4V7C6rcS3w2nvIhHN
hNdFQPabV0oarFRJ1emO7/5tAr3NVdKkMizZUZa89WOzzUao0IVysgN9nFVqdJfb
JFWTL4FIaJBH1JBQytt+QbaQuJEf01qKXddqxCCVDeGpyLubeYFGBdf9+rH5TNQB
bTn876b03l4J4sdCjSJ7DV8K+tcHT495RbUpMN0IBI6llUCyAHzt7tqLR7SlOQ6o
xO0qUywcjFPyJyU8NA0At6JF8JmMJGhg0aFDHCNnRAhclEPCa/RXrO2YTOt4nQIC
7JMY6PDB4iQhy2LsLnbQBJgVlE70fhx7r6W2vpMDY+AASuLmF9S1HX22+DAiKU+r
Mnit/dmWa7WVJa704+yqi3szK+K8Lqmpbi+ElfPmE6e0QKr9zZkMAe7CL5peOPoJ
lgtbKv9Xreu5Fjic6l8uZcoGVEczIGvMZ2UCDBud0UbtHEh5Vgyj436JRCXoQMiB
p1UfG3NHFSOpQ8XHdu3fnswnNzHOMmh64DnrEOygTCmlCne8Un7USXMaUOSjQ+QW
5MBZnL6cLBK6OoM8d37v+D0B357u1F6ly9U8ymQG2ooVYVv0IeEcQsJRXqECaUnL
sGei5I7lTNcfQ9sNg73mFGK+453JYCizphJEJRcfy7tUyGkrOp6lDBoKppeUrmdW
9TyXBZGPe1Nl4lTyj1TBcdsA1IbNtyeyC7fYG6haZ3WnRj3mq4bwPIaLnDdoVSZG
QBssTCVwLqKuHI3QSxonoowAUCE20ekaGDTKuWHYKfxj3CHyQH5slqX6rbjpI0Vo
3f7K2Oe2uHOFXgDUK/3d0JiUNlQ/9CSPa+VxjTkvadxQj+ipqjsxhBAdBPX0WQvN
9Ptg7HsbGSSl5gBJUuFi24tEhMRIUdyO07tBIZVgfhzZ1z8Wq/2IqM0gs1BOk7aR
eHQAb0pr3GCW9cdFAL9NWKlXEsE2HRVgAU2AhPJpidhT+BvvxkA2ENEPi2Cfq2sj
+kT0RD0zxavgvWQZETmNqTRRZJdVC5bhCkv2IXezGLSwNUNNjC9VcDi7xSI4iPdo
BdAV7e2O1u8a+iQIU9OMvsD3ciAO5lwls9KHqUu/drdTbHxfzzrYD8/H36ZnQnLf
ZBo1+RFq7/KBEumB8DptqqDD4BUCDBf/A87S+rgRuUpuIYRN9kV0cfW6tnDx9QGD
j1aAXWU1MMoBzu4J09cz7wZRZDyE8otxHU9HYEqybF481pniM/8PLuFjD8ttq/Zx
gUZei1/1UnZZxAyhjBz+/I/dfh7vfKGbmNLFYPdYeXLbyIRybh8nosnAHLDFkyt5
eVEtkmb+4IN4ba1/um/ORV10FX8ASu5s36Vz4N8gwOW9H4FX/P69QUY/Sj4vX0rB
tiMBchUk3iNJIuOPAbWU5wQaMOtEiI9skvrpKbBIzJR/i8cuxPF7B4lt9kpINnpU
TMrJx7Y+nTOeg36BTd0PmIINhIMKttwIgTHHxXw8LelCamr8hkljvurxafXNHVe6
fmYXIIjpG4hZGivp7GqXMPA3Z6brK3jFalzIjgvuHp3uRy3W+/iCrZAD9kZA/9lW
yOnQJ2C/q5ay1sSRswIGR1l0T+cepU4olg+d3Uqj62R1qoEGmhcRmiW2QZ3KFMSG
euG4x8hSwls3Hj+YNWDNXT7ProJlVChtkfG0hT+Lcq7NGWwhtLmV24tnOFcy4JpM
PH0yNJuAzbzWVOT3flgR6iPzMDUD9ajtJtCBNrgCnyPxz9FezDgF6QYAiwArH006
vguMlCIHrzKKk5y2FTarKTwsxea5QkrUZZeduUKKK/DGux1lC8ohtOA/rw2ACR17
Fug4fyV219eGwdXcyA74NSlIldakg1CGqK2tDYTxQGYOdKWPMcirwgjGWX2IsMgT
xOyGpqqi/kvM6hPd2d+FxBaKLH5JEnuVbdc+AZomA4o8AoUHQgPpYBwmiXeLTNhn
8LXOLXR8IRjXWpPAiMOG3bgClu2ygN/gN8GqpUaUR/nxQ9oAYS9cYuc/WHfwDjgO
3ViwsQnylxwfFIF0wVzQ06AnLtEPekidTQ6XrdJUrm6B3azAi0302OFZA+4d4Flw
RYQ7vKhM+vMLJy+PqfCpPtAKkcIBP5IgBUgY6EpsPi+R6EUqGdfadRVqDr3tD9MH
7hA3uM3NU0JnBBSpec9Wejr2TTMHyx8AV3j8j7bQZh3j3JArDdYDBdnKxKEkLA4X
rtup2I/eSnFST+bfBpQHpKXIf1UrWTYIGLpiMw3P39LvP3v7F4FtLDX7HgI08ULv
cZkLsl373Zo7xLiQpmpCLVjOIrhzsnM6O6G0t1joKOs4s4tkQQ4toxz72wsA5tqX
Z2WVg31g0ThHKO3CmzhieJ/MHANeEyWFh+iUV5KqyrKS75fkXHg4xtZxU7uY6y92
s/dFKtsOpZiU+55qLnLLjJmJy39j2u7a5Nkpcm9LUaaA/OjNallXLE206SIcYiGh
eD5BraEwIv7DwNtKRmCkS7H1Ow/KkyRy/RK/ms/e9yqG19gmR14DcjhqFlAs4cRl
P37POAPD7YU4qlxEJWFap+4AH9pjIIfSGU/Ui7GUJf3jnZwgc2+pIFMsWnFQ1F9Y
X9tUoI/3zonq5zc13gbQ9hhOTkLSt7CqDVNJS+q0wPK4DXkYDwWe/gOFEe8A1xLc
DAFj5JH9blXa9Y78QGrkqjp+hMZ2FxPHzv9TGYrpDGrJmPp5rIltQGOvq81LtErz
0ToIcWbCl1gUT5fo/i4BDwu+b/hwr1gphcv/Bi6mVzaoT9xhwmjoUEVVwoKudHpY
2H+Eajf1Wc3KSaxCr6QdG3fG0/Kzt/XfWR2E5WE3hg91SPRJDI8M3GDA+UpuvE0M
7MxYzs5GeEKtu+7Pnm28Ifk3pgJ0Njy8WLEUqZxDIzmLc6TihL93vAQJ4btSVm4H
6zjLFGjt3599vTcQfYMxbn1/yYghmBR3vCDimYK+EjXm1xFz/+G44bAV0RJFKbM8
ERFF6pdEC4X8L9900VQ+APP8M4DXaP1lrWKtIg9wxtihAb1PQ8dbm+qPRuqOozoX
sfh16krcFumz8UrKSO+OznEJTsGbat2jRgnjQjGflzmsrkk1MvSdHAVaWrXQwAdJ
V+6rQonu0qg+V6lhVQURJ86LeCpgEMCsnf3w/P6wj6ZoqnKSKa7NTbNYXp7p0e9N
N9X9fB4vTq4sJ8uK50gQlDX+eDWb3wTJKGAoXfwqg4l6sNnYVehJvO3oDJ9JiY78
FejU8arzL08DHwvwx9qBZoqEIIZRoEDkCnJmWjSdrDEirfrdDTCBV5xDUxUM8NOn
WkVU8BPMXYAx0KIM6mU/clR1pKfyinpggr3EeBugQcAf1++0zdDtL/2TWMF1uZIW
7GXUYpegBiTJyNY/YfD/x+o1uU3tOS5txycID8hUU7WXz1N+y41v8Xgl9qn5ou3X
nb1uAPuvUPz5dmW3xNvp+dXa4WtSYWx0481qBMdGHtlXOb7SnInauWy3CQMwF4C0
J/EsbQBEyXNUC9hWVVuFw+I8PXFqGgJm7GR9+h9iVydXIJpBTTh6UvdvL/3hE7Uo
sYFVX3xIriKZjbTl8IhcvJXTrn14/CcXs9dKkNQdlq5NKXa4gC/TTlfIhUnsDo9c
ee6gc26xMy992+xy5KICAI7idqGspKf6vUG2rwSbg6QDprLNfsiP2YjiKeJgsb3y
KjWwsPjmBdxDUenuHGZEXv4wa1RbtxprOR74L55knUog/pc31YBtCTnz25z0+qzj
fQFneMjLNLmHQMsg1n7dswEHGJnK4WiaqBLgtE1sjilFGUBxUoKtQVaCe4nrT+Fo
O85ve6v5KIycY8muq5E7c/SDniiaeHzCoC1sEFpD0HGma9JDqvph+yrPfACiES1p
E6ghMXcg8h1hvQbv/Vdfjrzgi/xYYLNeMGQ8OvPS36tOxI6dOD8a4zcOljqrSwOR
W8giw8Q1amIuchezE0dw0yuqPev6CGEUSOWhSYwL6+3UxPqan+5uxUO+BPObI1EC
1x/3OwMzKjcSqjEGUGFFhwgwXm1FLRfPd1iFs0zPTs+WSpFqdLmlZsfz13yRGRtz
cItVPCAq5uMKnPdRE62Fve3Hthy9oQ37QiOPkggTUSuIn9Xe/l6NMP9yeQ9zBIes
AHVGHCD/7J9m0sGKLS7xTnRMIJl7+yHPHssor3uLmuQpgH+X1ooV6MRnKPcbtgJp
q9Eo20VxGpJQveaP701+Jj+xgbMFsrCSoQTStHJ+aI3QaWqextMThZZtaEDP7+5v
Q7uH3wZzVV+xXtioToiCW3K9PMZhD2j4cuPGqTI3BAtt1yOfqLDVfCiZq4fCEnob
pFtPhUtu35Xon+CwaUK7iC/KbAK3xaJYUlSLbRNx4usSMw0OHs6HQAvFEIcE26g4
OxfJUNCm4vg2QF8dkDrDyBpzw+lEbRYGqAF1F3zcry4NXMw0RnpPZOqC68cCiF5b
lGZ8pl3if++G15v+PqRMwLwqY5VfIUotn/XonLvArxZdLQIL/IoMmPYiRWWOVjZ+
W3dT0TV71CfovwwpbbA3OKNZCyRh4jxX4w7rlmUVA+XQmWsC2cs8Ovph8D0SLjHT
I4u5M9++OA5uGgRARIvwE5kZ/4kDeIMRgKRsCpliKuco7dKRQPQhKibTnDOImxGO
zWlHfBLVnjTymO99LWP4/yJ0TkV40ZH7bomLdgl6zCRg26tiRo3Jd50pX0rfDMKB
wmKWMtKuYqczeOtBjeGhv8NKMlT3dYP+38d2HDPvlosMeZ7b6CwFIicszIluSReE
gjknwmU4sowZQvTCIofLMSfCwsz/yskLR6hzm3FU/8g+H79VyCjzVHYdcU8SfEFo
4T29v4/ERNEyg4hFEau72QayIhrohhqfXBc7La1++Ld/nO56LtrxQE6/0oKjkuwu
iCr5VVXBdrJgEy/L76TlUijENMdy/pHESsPEqKJ2MmjXag8vfyYDzcp4H4KyCSpr
KBnHnAJDkOZmckX7Sc9Mm1lb3OFKI4w9JXo/GJYDo6AR1FHo/oHxJjW6xcAGHlkz
kiCPLvdWOiY0xqKJmrwtw9VRAnExCVyjELrxrwnBk0xWLf1QbWYEqV+ujvzi710c
Y6FyslUeveY6NIuRrAIJ/zh0rcxIBdLn8qiMugyijFXT2rcM6Z2UEcvvw/LtzM0Q
kun3bokORONPZ2wAs1hZiH5fN8GqVvaGbD7e2Fu19+ENXkadUyb/nI2mYs7SyTe1
YRb19SZKrPk9x/7X+m+QmhkEV4lQwCkrBS2bvO1YbsMSm/YNSPteTIcKLUVp8nl7
DP4AY1PoeEPBHj+OnwDnV7PQC7F32Qili7Gc2b4V2agsrhfcS3q2U+UIleZUCAjj
JPaDWaJLmBZq5/HfZriK5x3eSXBc8NOEdKzky4jBeBcGegZQOKi2kYxk//SKeozR
1dtWV7tA1BnqNd4qcz7f11rKjKNJ38cSQraTXgAm26iiFiKawSOKgnPq1z5rG5rt
E6Uvyyqo3V1vSVwdXG+U1zpaKs8ALe8HTMtehLpef9KUWswEK89tzSm8VKjyRG0e
YD3nAt/HLGcl4ozJH9yp6JR0ebAU9s/3AzZ4hQWBnO0ZU4zLYi6QGJ65tKLb7yGa
Pb0LhubQwQAzbracks48RlngcoGk3TgcXROj8rcu2AsdHL8bEzyk1EJocEZb6tOm
iBa/DyMfz4EPnbNRbnJGcGTY1O7naTCLa1duhrGEn0GDqNM5/weJkHzlbw+AJWAl
49Nx7v1J8Ob0zltXQUkrrhAX1dQ/xvn45yFF73/dAgFrfcRiZ+jWTJb5Jdmvmfn6
2SthEEQt12umoWC4Q+NQXGVMceXVbNqhv1N/TF20WXFZhjBwe81oSpxIB9PnfM56
SVl3dGCxsZzSGcdL7jjVNxtdO5MFfpu1lxbjStORU5CRCkqvHItz/CEzgmOcLYsr
RWz0STC3XSIuPJ85kUwP2fXK5GH/oEj16qmgqqEwfQ24X8d1rvrTpAjzUDY1d/BD
cN0kyTl+Y6kbWzer4/cBnhy4d21BEqj5V/s9KGUtNiAV0e6hDfqfvLwJvH/HdfRB
JiPtkSPKi7W/hIx4nO2TxgnNbDNyDo+l6nXoVoHMa2oEQU8lTlCxMb2BH1zgEYRb
qZIB2zEnel5PPj4WxV0in9rtxrM6di4uyfSPqV5j14tAfgP/RH05wgiYQJy1TWa6
m1l3CFAMuBYekPrAXcxP70t+DfL0BMUGhwx2MI+CMuk5nBGypFovN7X0VZ78yNDc
tjJKcww/ju5uJUpqwUcxujhpkaJHCuqPTDeA9BeRvRViv+onrL5voNxu4+XwirgO
Wdd/e4DwZ1uKQHTgE30WNvbKTUq9pYCvBZuLzrx4MENur/taZxo/CtdBNFFbN78j
3LmWAlsO2/HmmSYD8iMYScz2vTmpRLMEkZE5MPBgrD1g7gOunY5GJzUASyUHxOqW
zGiCu2ZNG7rOMEjjJOXTlV1mnWvCPRT8JP7GpDHejQVqPZ6DD7w/K03dBnQOusWM
/hSmWt6AO4pPeK5BJo3Vas66pPA7mWG23rf8yb4uuAZsv5qW1Lx7xJtC+T3tQGh1
C+/QqMpiCIeQmr/98PYx0tN5IFgu1mV4KRT13GSkLSuHh+qFgz/yQc+LtGKr/2pV
ylUxtU+v40ej1KlD/Ul45JAqGnsIxtrd/qvvQEO86dbKjJ/iYPSRqfD7jTQJnkz1
uMr4SNtICaO75rtWXb0AYdrP0Nkr+qmTA9bdgNBEt2umJrywaDLVicHDvITThhOa
f9kr+N0JIUjbtx/JZaw3IDy6j/D9hO6vhLXS8W5PHmMHlyQ+z+8qcQpvelRDOQ80
wDapiKoSQtWxsYRPIGpjZegkyU2Aj2RC9cD2nGklsPpCBkEISh2yZV4czgmSy2sZ
k54I4n/6GcJ9+NpnsJDCjFSdwg2GJ3IudJJXBLblYkGjLgYQXIxGqjRnrd5zDfV+
ssLY7qJI4fZgCbCmeN72EQg5owkVb9p6ebULCzyXxWSDjQ+pTwWYWuHzyBPfmtKG
WRIfmE5vmd/QZcCDoTNsJzhlmkN1Dr7yQrZv42Xk2MH6bxASsx8KpjcbDMY6zY3l
5gGiAtMayGsQqcpmu50whS9Oh4fHrtMYngATsxL8FVJ+PKnCOFC40O4JdspFrstJ
4EZ3099C6BERagKkW4pZemwElr9QAv6hoxTv5JQnAXqEFHn0XhL0uvWETSTtZX/O
4RY6S2o0pSRc9eXhMVY/XZbqNUpn4GNOoxanT67LBq76mvC2P3rHKJFxb+S1yOyH
rI7pw3CoDcCETxrb6VjrAGaOa2rJ6yvIrCCH5ekmfvguV4cYqca17SoF+qdc6mAl
HKIdoWAFdRT8/EiPPezmb02l3hPJa6iLYhcMgT5fpFOH1t1qfzXByjEPJJsZvhBC
EBF5WwJGf3XgOPHvsu+6/cerdEzSSNwiOFWyhLv4N6iqEladm9VjPOS/05heBhDq
NRZ1PTYgMyZJhrUL7H9bK/IgDx3qgdIWYQVHRp6DeT72dkwlmEDJx4tlj9IljT3D
U01ILkR8RhSPHd3dmrCsCrJZqID2i+O0POfuvfngcLReYRcXCiJ9hUt0WHfMQif3
5tFLwtWJd4oADKR5Qvle2rOHBUy8Grns++I7IYv8TqQUCTlQJ4ZxpmO+S5JxrLmn
kvgCb8oVyUgeM8lb09MRBOn5y1LQ9iedoRFNKGbzMYsXYFElV7S7UNcYpFbg8n8+
O+X0aoHqSyCCttMcHcJwVLBo8W31EfwvltYU73yj5eJ1VyEta3zzcQ4T/JqttVER
/EBTMtUaVwWGw2ik6c5RvO+ZXL7+5GPA+b4IEoDoAlXE6igyW1uHQZJNlk/Hm+Tm
UAmBhqUmzxTfSMXh6B/C8erz2OES4PgIbcAv/QVLaiyVq2xPp2Duz5NefhrOXtQW
UBxM/V2FaEexFCuOnus2kuekU/KeABOYj+3a4FwAtn6ZhgqiD2l56Q/LLRTcs/8T
u996m9DwAyNMwnFtI0D40RryDiKk0FdyZTJHLNEh7igZ+Ob6AYfAfKVnPJIfR9gd
9aSQ6hr2puZCU9KbmdOdTZeXnpiL80l1nO8O3LzdHjKaOpSUBNlBNmxhyfcTvahx
ge6j8YAj3TZdI+G0MtUwZCcOLAlBQJ0WGPcmBHwlPV+Ao2FBnxb3led8LJq8sQBX
yfbXtjpQi0xMeEaBGuxPRGNFKW5bA8U1YT22tZVuqOn1XNfL/CQwNOJKL1vYKBwE
9viXQj/77aOQNyshAMatzYa1F/XRE8UOXSnhbKwq0feHjQe6eSo3lhO+Qmdd42/V
rvdSm2h9ZETnCitIOIjaTINdag8bPM5dVS2Sgn1rc+SfXN37+dFfUm5lc6YpuAWJ
K+DiWkIA9ZFPSEW1/66B8jGDfkS04EePIGEAgvkpAVgN/+vrlFUrvOAElgZk2VlP
qhFvrbezjiRJmN89HZ4S0+bjlTj0DMMcPBzCXr+Mu8zQ+lMYAVWExxQk2Umcsax+
qzoznIj48KDg7Mzwiw4V/Hq1tD7Iw02UX54aQ5LH9FnCiAb62P/jITBcZnoh8ovv
EWNLmxiFFWFsLkGAY+i0xglXYQMfusqs3GhML6hm1c6vzTonGn9h3holKd476XH4
wmLf9vHd6k5DjIKHDKdk6Ska/RzucmJl3/J+4D/to+zrwVXaD0iFaih73obMVXpC
ufkDlbzi2nLXgFeoqLkA2CWaAZDkvvzdmczSCdHum9aQEHzggSmRRHv9Q7TLid7Y
eRBmKxRvYQO9h/9nc8sClmPbV8S6oPSNxokyorYAMQD4Z/jeAty+1JVtPOfirw2Z
EXaGghMIw0osa9JPUKAaGBA0IOmZJKWDVeQTJQE9rsSmfn/BcQaOEHAmny/Mzt6j
LHE1H7N4NYDJv3fo8gT5w7jqS6FUsmITjfEoWU4U74/xiLQYhlhiBWKO508wg2qC
EFPn/emWS0PPmqycpCk+xpVK21FCt7iQ1Z9Hm7NDjF5UxjdWZTLSQw3PFU8eQt4+
Rji/ME474bk/lK7U+q6Kkz+jUGtCMcE5+tHfqeHrGiQ+Ff2tSogx8MnnlU+JElfO
/TTMg5J/ZqssyquiMtwjUXBSc3IFhdRuJz8piugBcRsy0Buwip8CvOo7L/MVXyaj
iQDGoI+OpqWmYpnBiJ9oq+pv+IBSso89ZXjkpcqIhJWDgoea2Ucfm8dCqOFcznwS
rjtcXjql/e6uhADZdsFdTSfBiXKs+TCZtJVAzzzlt37O4yp5K/QFEyjMnCsrksD7
tD3VE8SE60LtuTvhjZN2Tdn6Qt9QGO0aPOL2pjSx7ks0DRRL42IFhcwxrpC55Qpw
53NIcr394oEfB7ygxiIOSOHKsdPtSouC/B8GKOWCsEQfKGDcF6dow41INOvUO/fi
A3jhz73Eg9AzJz71rbGCRKJuhlbbTx4ADFORlv7bV5VTcNufGhPuZNdwE3S+6YLL
ewFKojqBzumBTzDrYZKfguHu27UXHhtdCDql9t580pyNGttSO1yub+2nX//dZte9
5QNieLlHajInhR6f6Dzn45hL+8d/5DOn7XBSqPGLSijc159/fyAgDX9BUxQL68Ru
WuWkbCijOm6cmu8fIL/F5bGIckEnPyfNJtoVUc85qjCC3QVRsN8MBte6b/VfFWA5
O2V8kWkMuZPaU6jCHttIG2yjEU1mgM6sDa3pzTt6dt0X8X+hnN+dMBIIaBlF0IrU
pWBbxSopG4OUSRb0cCZrnX5CTG5aSKNElCg/Kq3ms1wfkUzBh91U5/6ofZuCd2fh
y51EdKz57qDiYA/66eNOs5GEKOAPq82Fqx5RtHNdzp43CgoMziEZjkuWYj9Uv71J
iWslKPINeIudQq+MqpI5hJ22Qb2XFwy2he4aVUlEIro3m7vx/2IYjnU+V5tKZwuW
bX+DxZL5/f3mFSZTw7KWRrfeUMl4i0FilBCuSMKTdWVArQ1VbofBfOBZKYxExJSb
T8ea8OTY1GZrnZFV4Z0ZppuF1BUy2DVS33efefCXSsFTcfGLmmLJiv7Gt6dGQIrt
1309zYoFSZnf6LF0ZVYQLXD+rEejriaB1OMscAunGO3ngPpKHQ48AUhpx8ceUEwE
qCM54Z23LDQwLZp4kxCZgXuZrekZ7p34x7lhJzsoMFVGZ8a0Ailspzf9yqRXOMjX
JzhV8+3wAFHGKxxSaAvhWRqqYsH142yeIpyy3TlF7RRGl4ghA5gcNilLYhzlcfgX
EVHCzvv63Cp1pfsYELmPWWWCE685HKpDeECic0rE7BFhpi+0OdP8Hn5o0BIBFi4N
NpU4I2MWBW/XzcYrVZ5tDas7Eygmb+GAi6RAohMf80cifn2KnV2R22s042GaJ20G
EoYMMJ0EMaGZqSTF10B9IDbqkyYt9zq0arIN0StbWy1+DhTptxuHfOATJpRVLBGS
Z2BgcB/lYCF9U5SKo+yfOxEmt8f3esqqmk+xBgglrtM3sBOSVJtHpRzr5n4cPMch
09pwWGVsBFGZqZiNITJKMGnNenr5XaFUzoyfEmeCSU6w/4ISw+XPoO1M4jmHuQso
6MO5G3Im1gPJdETBQ4QTvF9sFccLHrXG/8l4HTpRrFcpBEUp9dwIOu+5ziaoj/2E
oAwbClkPbKw+ntRUUwSR7xeqDyzoHLslguBLyS4kEIV+PElMluGvxF8YIL6MPC5g
XTBXnWZz9wA00eWq5FWj+rYMSTQVw/W6HQCQgFQJD1rPBcnC2WuE9d8CwoSkw2iq
+W1iHx/T/3PL6iqA/chbcEeulWkRLnok6oV7EgNPt00trI+pscESHFyKABpoLDiE
pAZUAFtaXgHQql8oEauK/j+8y71FXSwAmiMs+iCLAIlk9ZA+G7t34ZTIyAqV6aNh
ZhaPBnNMEsJEpT8pBAKMyvRtSfGLijEwq25jkXJdkt0fQsRvoM4cDIzUX9wdZBsx
+0UzFS1bXGAD/nT8UbDPpuBtqQPsZIHcI9zC6c1zRd023AeJtsNML6KQz8QFFEBq
lLCenoKtn0Inoux8OrP9+9OYFPWbfE5816B95AJNuBRbdy7IKBMe5jWjzpbqAQmV
zkXrDtdcFfrriqO0OiPnTU2jn6t8JMZ/zWx+/ScSPJxhx2dxiNhkhWoyLeRhBJXw
qyyJO3GIZzeAiz/OwriG76DJntUQVRgM0AXH0luZFfiu8FHClRoxN0qmORWCNfHv
SyPKY071W+teq8WwzKUjZrudctxoNg1S8jbNRkqm9TtpBn8Ahn/YDWbJ6gulGfOi
Uw0glwSuhd1yzIH7yEzKymbSFOXWP3b4F0lubu292hXC6aY/4JUIStIRdUfF9aT4
M1p2aYq2bk+5lOrU7KvsSWcW72titr174cXat2kXk2cRdwaXP5xXvsHpwmkHyK3N
EIOlkcqltjIG9N72GsZb2oacLwms9igD1oATKso2MFU/hgB7Ssf31syJfYqD9u11
vyKDb9xeMgoIlaqSYZ7vbwOM74YPky8OV0wad1A54Yr2QkwRxCc3xU/UfOV/POVd
Hmm1LXDDvDLBcPgwv3BNfmmKbFhNSlmxy3igSmi8nAAZHywxIvF74rCcuUIGSGIx
5vL0ZWp+YM4J/cWc3LrgMZa2GMbzj9N4NtYRqCvZbOnezJyEXkbhWDoL/i23Ssjd
9RT/kuFiAjmft0ybxMJNH4H8O2jRIN09CgXkBO+6XqG5Mvhyv4+Ot9uiQho9Mp4a
QHPmcC0xQMpFdf+xkrm5xIR1jayIFyRz0x0TqDCr4P4dqJEH6hspFrzivt74vygJ
F6Twk+GZZztNQvtSh13sh+FndTeX9FMqLV3wHu9HoytYjwPCnYnMfjupUAeyVBE6
9rcFS5j2KKA06IBFIKzVD79HnqKd/EUfrZdjbamnGNB7BtdJPm0jUfOJH0SCXl0e
prgVOS/a47brB8xY5mRggQwULfWwmLfdnNa2F0Ek16rWChJxjcjl+GXRHCT327AJ
80U3Z25QI+o6vn/PDPkxmODXifYxQmtrx54T6RlScfjoZyixi7+b6XdrPd1sHjoO
Q4ow7Kkn3QKbnGpkI56Ul72ThQ4lNKcPnL9YbPj68m5YqzpXrY9uwYR+jeQbsUQZ
M6jh79lpvI1fr8zNV4jTRusErEuVaKupiiSrHIvCQo0OSt2Tpzn01fBmUIi2Dq5s
3Av72cNFXS/7fLHBk/mGyjyWIgBRyhBMgrZWWsn/b/PJ2dG/QT/yCgzvh+mg1k+3
s6Un9K8RIlv9miXmDgOqZkLOM7l1CrBdwUSnCGJ79TAQ2/86zHJNLCwPHoyaxO+z
8GeZyEotnlRomwZo4YemMSlDS1EI564PBYdbqAyZUkaHkMwX/fP8Oydj9fREsOMb
4jCDH7Bs2QibJq33+k3eWZHZIn8/eRTsVywUTi90boeSS2N9UU9AmwZWz9zVmVZm
qCR/ahd5Rgr5mZ5ZpaBEQomP/hguZEDTwOWtmvPs04i9exfhkyNXqboC58yRr9/i
N+/0IEyJcFIr54a6q/34WwFnvjGq+YhnyVkPLTB47T1AFzgDE0+wl3eqmB11I+cn
6uXESFlHg8+vDvbUVYbc/jnJR5KDBbbiUmSOVeFjVmyPd3e+90WRLOWdAMoxkUiJ
CPttTd/T5nct9t+lsGjGWwtJ7VH0NslvZ7tbuDHPWc/eZjw4G/jqQJojLGZ+yV48
r/chR0XbRWrI+KryvyUhwUXv9lVpozu3lLGtOLUZX4j9MZe2ni28FVpoOX3FHtU1
bCAikx7gOqyKo3fb78eKR7JfwphUyJrL7bXOWk9n4sLPdHUB0B63wehbv8cYdUpP
f12EJjDdeiViw02TxEq2Yj8MHxMg6il05Z1DlPsnIcsjdWkoWnxjmW8NF+gfbHzA
sGdckVe0Q06Xn494pCA0pfphup+yCs1BspGuYQinEKbI7VwfdvfUHmPrOvwHzMC+
3N/DAlJzPFgtSKAapbhVvmZAzn3n94n3xdF4XxpIw4K56/KCr6ZfF3JPv+bnSx65
PX3nJePWNGU1WqTnafr0ciKCpfxzdLbp2KN+TttSme8xcMbb4uEVf4rpsjaxCoFX
yxgZrA0JVBmNZNRxAW5/AQY8US2aZ1IoQdGOx7WzO1ynLildvm0vjsG7/BZoVd1t
f6vQO1iCh4yutajp7D5QsebMxZ+oSxdY+vDJSvK3PXXsxcMSsPBXFLgSJA470WGc
gGHj6bIWGwK3q+hN23MwauRp4PIrIg8PR0/9DtoR1hP4VXMO+xqPafVchN3jijif
a8iOYQbxfQ8axcouQaP9cDPp0mjXp/5D/plp2THTlxI7CdNMhPoLvfDxcN/fdAcE
uGSL7lopCAQ7thCP+gDAwR0QkxhNR+wtWM4UeoHtuYXVPqipK8zdI4Fo/Q2k71FA
b0ywH/DpJqpa3CR2Rthirxj1BfP6e6DaKqkCVJ7+Krl5vPUa8/F754sI0zow9dlt
/J3wTvPSYMZH4KuZXtevIoHjToXwQsQXayCMaD6JIEpmuPMVe39Vp/AHsUk24Bue
eNXmF6Anv5BeQMFhSF4+uSQArMuHily/Hr/DJOMWpnGCp7vIPc+M+TQbelQqqGD+
C+TcIYrS3MUC6zTsPf2L/roEUq+l5H/qamDpTBI3gy2KRv6wXp8BWdFpcAEmp0Xq
ddo6bjCqDyoxQ0PfaP6810UXHka0d5xlfNLumKb4bkrd+K7pTK2mJFBUQWkeBSkN
vbSmKEev4gmJo0lhuOLvrMECEIiT/RXVE2DuE2LsMEdyV3IVfX+Q6znk5UTk8VMW
M1rlHL/ObVnbKDtNb+aSvPkzQsV9rk4boEDkt/gkMfhW6VMHXKtKCDAnPqdQgAQB
trqpgOU5ZvR1o/KpmXnaff17wBAx/tN4zkgZZ4N2biKC64+NAxzN6JWikfZs1uCc
DvuA9E1sYl4O4qNHecPCoVIEfH9sy8kduLB4GJqoXh/xX15Tx/DrBhE6t4KW2Xsn
ywzOwPEiOBalcUwmvxJRz5lXH4GBTBrh73Bg3o/73wgh1PJoc+HqzrBuGDOhOYIj
+reRwsFVaLZ3tySkb7lgSualv26kyZ1tV7JWjgH6l/5LOxAcVntA3na8a8cTlloN
sjpXK5B/b7tGCoTKmq4JVOlFddy0Ky4ZpsYCl1F/vZ7IHFvBUZb+ktc+2wXCyokT
Zj9AEzamzjutjrNzlK1lvg6j2vJA37zK9GAg44h70hVSG1JwIkSg9+LZ2XiOutFX
MXbokZ7xfXttiz7goA5JlQ35FSZfDzSdUgYRX5f5XERbkxGEZfDjjIEhMAmODxNU
0tse/I5vv/B2lZ5kTwQkhBwkpAxvYQ2DsSlAV6Kwo/CJUBTDKD1MeTZ9CgOOMTGn
rrCUHtCRmFGRA7fpThhM0Kpvp0B/nmFpqsVGDSgZD733Se4U7BVR3CkZuVaCtQVK
yTMkPeCwjZbAT7zEUqNOZXJPVTpPj2Dj4PcvnBB1pqmrl6FDXeENeMhdu2EHaHsE
jemNllXaWsn1BjqVhXCGwVpdfvzTdtdghJzaWTzIsncf8Eni6aOENtQI9FOQebks
/FyPrc1DiVA+gA7oquYrdYxhVd5Euhyvgz5hJbUP7VDzNKrR3kYQ7uw5fpt0yFQ0
U6uw/3R04yfdYFQ0/gbmBPgDI6Lka72mA6gL28061AjwVof9q2+VWzi+ih3Y1M7h
t5zjcNMGl0YPNZVNUg1TzFjw1H9vQH76FomnG046f8W0cMd7DmA8yc7CyCMVvho9
xnCIJx10T29XqdoaKXP22umznCkusnVoTuq4Ri1LxvI8+yKi8gqIB17MDCqbh2jU
Rm8wnOnc5HQXkyB2Wk8I7nNI19tZpwBhvj1Op62FphRO0bOs5w0ydNZwrwGN0AWB
pLMzcokfiJwSC8hLP1ZbXqLES10zETMNXJfYta3ku+g+vopGZCs/WY2fFgBhMf/J
WjFNhEAhg0Hk1mF+/rs7pPQE39DLYwj2F7BBI7iu/UyiYNLkA1t/bBNt8TwHhr33
lSGSbCgLaHsZDvoVgCM7I5ctXXqE9f43kJamrXKRwhBYqaasAKN5NZiWsnk3hRVS
/oMdu+itWlz+bEP3bgKJGKCTOko36PdUEYaxiEovNCjBnR4TzsIN8Jv0CIj/67LM
7BporxfU3VYvVHVAUbJAJa2Zvb85wYy/5/ImwPyzlWV/BQSkmD3Xac+Y/2zeVG/t
2oAJdPMEczDJfUnVCqlSQphGo6dpv5dw5f5Pe7DTmFcFakAniyNv3maBvfjUGiaV
pklONEwNDnHez9fFZRaPVYtLT/I/ahqDD5zysNGe+p5I9JBa/w65nX3/m9vj3oBe
G4t73cfVli8JYZo3tyBDFW2tVPyK374Y//L3Mcl/kBk81LypG8TxkU89uGvjRiQ8
/ZvIlphCOk0E9IBB9K47FFDbLKWyFkBgYLIaHJu/tbXhNHX1gL7LO0ogryiFEpce
WpgbrfH5ybqGAuB0V5+hGsARic0HB/Gbj5XcskH86QP3vHuB+es/eCJasOykjnjm
r4yToXfgHSwCK2RI+eERwh9EkzO364zdD03ildeaCsuTIGP7i8lwsNGPgqF0c6XN
NXl55GbA+QDQulcVXh4//nkMltsA04eHviQThX8Ma21gaMbCkoc1T+vMOjgxp5WA
WOZKT4X8NGx/JgLUqx2e2qhvo1ae6ymdVAZJVrIZ32rGmxucuhjhMfI6dv0SsGng
WQtQg0xYgdss6bCrnr7vgMB3UDRPbRQ3dFTzbeqcoQM+Q/xx005WjIOS5qVzGbKv
W56euQJ8X2Jgx8+8g6y+Yo9wakgpHCL5K5Im3p/3ZH2UTIL5EqghPyu449eh+7QA
36kC7Ki/0p5DSZZubvBM6PU4KuodOkUzlxgNlcDKg0W5n6CvNQgpxyvHXEilO+V7
HSl/UjSkH3TN/Jr60VVuph20dawbDimPF7K4MyRa1rXe+OlAQF3DLlWcGkJlgFCX
AMeh/H6Smyi6rcxmTJyT3hKPqAuylqTTxkggh4kuGv7anaEYjJkq6yiRXs6u1xag
47O21tfp+VQGweER+SaBXDuJkfA9nHUkeEkNgCkh70wasJ8JT+sKQ6DZOcVnlwl5
A57sKB+pFjr+BwxJ4kjkXuBegYqCUvRwSWVSuaei8S6Wl0sW3Ky9QOBT8ViZPSwK
p3pW0GZEQIndSOJzH57WruBEHKttqrbW1kykh0/GMPkEE8mIHiTy4KyS5CVyHiqR
jYtwvSlWM1dNw4YOPiCPH5iF4LMNHZjBuK+by2UC4hCVgf37Yry55Qvnlp503R1l
Cev2Dzfkl47CEk7z/riYP8n2SvGCVO/PacMdNGqU6FT4PihpYkYFrP401XAUUWWc
36/va+4lIsY+jyoxjTWiTGZ2dHPpsLW3XCEKGhrsMjPsoYYWMEOvACSD45fPcqXW
kTtgYiQbTZkYgTm7avjomypgkYkJQM/x+iei84oxwTi6HXs8Co3iIVMQN83Oppzk
djzhGxyEiUMiBFyzsOVKiyi/X5VoarGqQlphLdLCI2Z3EjQzsQ6UsBK4ehkeYbhj
SpplUHkD9FYh4gy+Hsyh5NfKIbzGEo23+CLyUdO8G2R6mYcu0VaDYHROokH1qju4
jiHG1e40tQ5cM5nKhJOFh6wY3G4aah04/0Gus+JjvcaKWkBryo42P6h3CJ3qgBZB
DyCkeVy5voBiCwhRYfUpvLTMo6bzVqdMwxNXRuSIqkNIlL2VonR3nxg6qF9crRlz
KPILCYXVXVAVlhiu70pN5t3+IdIa02YQlMz1ewTIvxKrP8rU3EvCThUwjshheEDl
6IHWJf2qcvqVWfws4neo5kUHKMR3sUWon0P4iDO8nAGCzgbASFUUYloWb20nfD/b
j+lMe9TiscKRPMruOK/FugiQIQRJeMkmxeS8lq1DNe4ifoTQOv7aYje/icPncXHw
/R3GfqqUXplVV1doPqJtxtgetVdumsR0y+9boQsyW45qJmNpf9HISygPel+14rcy
gdklDZPXPgJ8jUPcBTD6+HWVgLLODHrXvqbAPgpQFBoeKjjxK/IKSgWeZBKSRxrA
cS/ttVWRfaAJ2K9KDHSMJNc+f+Zn/kVB/+dpd3gnU7w5mWzz0mzlfjHwVnHUcPQg
+nNX2eVKeC6YBGmReIk5Gqe9L55nScrKspTmbOw3/qiyBqrvUqq96W9r3YOBC5L4
jBoSr7TwZYvGmOR6rLo+Op9S8iCN0uTQSWWHwI+r4HxXsWrsWDUy8HzBfwsSfNWA
21et2CoU8lH3mc4whwXY/d2Wpu1NrqrBdyuwWY25gsCRd6BSEC3eZhVCjZdfBP5N
HlPMaieiLJsdWLoHk6aEQC7vwWQ/9oLExEXONaohAdKA6eBgKPHgjv/Z7o3ECJDO
PiEA5e2EXZU0dFzYgplaeTZvIIGKopum4DvCprojASeoFvUOXi23fEjZnYAaJ2o7
50MX6cMFGdbhe4nGJTVySatUFL53vbD1mCTGY74PJ9fJVgH6UpYfo1Jb2qsnZVSk
ve89L+ZI2FBS1Dc57d2pQ2T2TdCBJxsJ+PCxYgyBInEZcppf2wxkCwR9XFDUTeAy
LCbktP8Eoqr94SsiuiFyo6g8e60B9lis8QGRRrVLUecqN3RgrfTLdTXyIBCCPO11
HM3Noc4R5hfkOYw9568O6AnLSlwU1JybY4ZGDhQznyYrZpf+64GuwqFn0P+xubWN
kBzbNVKM5UYCLaXBXNBbt2gWjyoNIBcTNke+SwxDIA0tDQDaya+w92SpfufW0fEv
TlGWI34kN44KajfQBncM5T7BY/ga2MhGHHJzkmsfPwY/s5gq6sxRor3J5OguAUJ+
n+uysyMv3qKCfKCI3z95K+1PSp5sWRDOXbpWnPe3AwbcgUxfn/E6I6dDeYvDOjck
kg7EumnYqerxfvS/SV6PY+UyIV2XS6kKuNlGMcEWpQoMryJ8hWIX4crrw9mtQfkg
+b0aRK4cf0EIK+blwqaZeEq2IqL3KbGpAiEKJTrhztbpH3nDZuVbcJmCASfQAow0
7MuRGNvJBql+uNIQolETF3vCT/FLlOxMuFfTtVq3IU91Bwsx6KZH2Kygtkid54vI
kY+XZycMH0czE0xf0cw/PIw9bcWzgneGu0TybrQ4U0dQ91ajk/cUuQQEICCtljMR
5zI9591myoqyuCatx2mr5MAZdx/TD/mmOyqSQhjqn2uPGDqPlUnxwiRNyTYZgdCk
bHVs05Dd5au/7gYlyNYgWmkaOmOZhuozYVWPy9VlLdME3I4u7Dm5MMMII6hk12sI
yrJF4xuSnbWL/PSt0QTKdxnNTWFL8QQs7WrFQUoJMfoNv4RcT6SrRaMHeqg/7d0w
R/W41lm7sY5E0XsJ4EE+Npx4fa+4IVl36BSaqVy98yck0KDyWJTeN0pyTqYOIqji
C3DPzo2DLh0Wn5zJNmVWO5QW0lLCC0q3J8X5R75foUSphA1KNxdPXqgsDHdyPPd0
2igciR1p0lr/pEovI0HpmcA12e/HmxuFmbkV29ANbZF8eofcvTLwQRKD0psmXaEW
QrTDR6W6YQBORDdBQXF39skh1i5eRfubw/r8W+UrGd+zObTv/Quq+GRkCvKTgAxL
zFrUUlSdDQL9EUvfTsbzxFqgcFbBdElpOw5g5pyaDpP6UUtLeMbe3KLlDQyOzy/4
wb26+7XSYqu/uUfZxCWubINXhT02rEenRpJub6tdfN3T4ZUBCI5aF5Tl3HCPHeo2
b2I4Gw9xQ6TrSVPKpt+GnHoKOpl+YGDw1u5M+Qqrlzeyfd5nZOhni5DIIIGYvAeB
zf1g4YAT6YiQlmfkVMCHA+30vORe2y5DP/BTqdIe00x09XyVhr8GIUj63QqIuN2+
eI3FO3dAqMICJMlCF3e8m6CeqmJremRoPoY+k77YaTfOtZ6GRe5vuehDyrJHbwpL
aNGUCAgfjw/OF5iMsiMXaOqyhFed2U7MlWdcPMJpTLYyqj/2Ydc7fL1lJ84amNy3
zE9sYJHKMrFZEucLn9SDcdf1ngTYtiUbsKTzzDiFiaYV5fD+fTPq75F0uoWflTKc
OYYiREDnUdaCi8BwMBg1M5nuEo0gxcVNzTRcu7cYOOXdxaaXziKCeTzcKDB1TXH1
RY5lTAWyk9giMem06MKH7KO1/Nf+IQiUPCug9KjnW91vDZiavr2aVkR12CGdd3xz
QMxcpP7o6CYLkwwZ9opFbd4vKvUTnQK/Q/cdXwo7CUf28AqpSL3Al90YEFA7AyaI
wgTHTYEKL1cbmHuafMKbDTFTkcsMuxHfFFEpzZANhkGlRdalULv+9Wamy0Ft8aUl
DjdxtvspELH/jjBa7uk2RIFQyMgIy0D3WDKY5phhJFbqQpjCI70fsO1IPYLOJxzK
JHagTNjFInlEaq96E8XR4L3bq32WOzT6BPHhSv3DOfi8Vtrhl/lqn6+sWlZruS8m
I83GJfZKKLVLwQsaKbTPH30cOTc9+9yDWzqdBvyXOjj8CKE7tu4y2Z2ke+v5tVj1
0qBXP2xb6GK42NTzjo27nXlJTLewf7uOZ54bAoJ1/uX+a4YbUw2sFcneAjrXbkY2
FP9YsBbHorlDU/3Ox1v2UIBAPTciC9BbhP5T3X1KKM9OwJr96V4ZiolOxJlGyOOz
JlOSRO/eLMb3w3/ih3nbN74P0ZM0ccxrwq7H0Zq5VR/77Hf6gqE9y4037JYAg4bD
dLN0X2mzn8ew4UQw8DjJz40/RxEWSKqM1+5uK0SPxOsE1c8Lq7oN1BFcbHhYFhri
Jq2CqfZ1pHXMenqDhQ3F4oKzrBApNIvkqOvYfkqQmimIfn4F7XLNEFfVO387PR+C
UNILDu0R8FNBjxNtwQdJRz2zc66O9NIzTccxWj0zLliZMYilsXFc44gXGmi9Mz/W
XqFbGOzGsExG5pwh5ryTL63Vx/nbFEIrmyxROUZESijF+KI38hw3LQp8wjVNXTN8
bpt8fiVMwI5tM+VvfkUbTuhIZTKit+ZqR5G5NaVtiF/dLbcMsOJvtj2OF5QwZwC1
vTqJDh3R54nVXbjrtOO4dIK85nKWzBvXP9XszBTUzthovXrtSvZvuiCw4jyLjIpW
ntduw1zT7FrUZC1AvUgn5TRivlIkPn4UUoS1vkgn4dJrPsP7v7JN0jy5/t2s8KU3
NXLi2hDSnHmM6EPy/g6l1+g+uCF0cUqjrdw0ltGAR8lAKXVGB6VObpEj+wLp66zQ
Wpxu/ZpouA4i/SffN3ftN0Y09vNayKTS3kVEgQsWv0Z8RIhb/n3brfM4ep1JErZI
pOjSK5ocDQCY0rrf2MTShkZSWg44v5BbhB2LSky2f2cN26gyWNcbY0NdckVqEtk+
SRsWGGgO/VUkLmlIODzQogTJdT0XVvbqu4Xq3zx/xXtd+z8XdOfQL5sFaQBJd/1O
1sNTeZqDHj/H0yxTgCL6KdRWzp9EgagLayws5B/Je/adWfVt0a0wRtE8rjmhwG5G
tl01Lt7y7iGXbSeUba2ekkLcCuSSqdgdwIWS0gWc7alZoEV65XBxe/QR39iNoWOZ
IO47HT9nX6YxDXDfKokEoKp2G+kjVzPzLYylT40yeOPZyx3huMMPESdMMXOwJ9r9
acwwNSKBNVlIUJ4fnu8aSoljdhqFu96hl5/+nViqSl2hh0Y6F6mEOiCgnPJKwe1z
QIVc62Y8CJoLLDVbBquXuIugEj6JZca4ESbQCipD5avIY4K2hKwzH4/XtDNdVjjj
qwjc7jJOi3f9Z6CDILnUQHp0DEz1xzDIjIHyu5wFpvNz1TCbjpRNOPjSmHkwocX5
XZK06PV3fSHPBnCKLypMUlimCv1oiiwnDAQSIeK2VptxFwLQ6sj25UKCHSrvFTcJ
YTEwJy1YOx18BjktCy+x5V6hJj6MUkb1YkBTar/foMpU9rs+JBdBvTNvHCBTgU6y
3Lckkbrs4DwaQ6GsQOKXzuplpCGCswEcUdv4GCDCg4gD4O91of2/Y/1CMKLHX5I9
PQ8hza6ULgSTpQJeKkNH3qnol3SegEg87ANHw+pPaiubkm/uAsmh7foe6l0LgCsU
fhGr2d7dxuIGf5DEYXje3BL+INdsY5H5hiLuVdVVOi01lSZLC9pe1h3rJoSobvxx
0uv2p7jftUdT6f6cV5a88l8FaJhI7FqgpN6tTS3giNqewTTfxdfFaFbPKvv17pdh
Eg45xVxXB36sk2tKftqWPd/b3c3mMcgsVfrI/5gnVUHaThj/x9xdwflzCiu1NUvw
hjsdlDc0CH2TWxNuiqfLbsitCZOoFvDTZom5V54YsFBxRY4TOAZGL16L+fvIZJZh
O58To4KMHYO5GK5ptb9cLPK2SsPtDIQrXTN9PM/X68FtEzYtIYROMZtFvlajftOe
iHrxsqG1miRdLdl/hLUz6o0QagfDTaGNo4rgTPgardBW8xTgM1Eif9pb41/RFTCU
pCOTFnsnoiaaC1ZSHG5wxsp7w6x7idv2gYbOY7KT8a8R1muu0KTxSvmhQmi4I3Do
IyQf6AfS6PbDs6cChdFP0VtfK6iJ4XYFfdPB9r2SacbnXRX/c1RMbxEOVmMvH9AX
aSdyt1G3eQHgtJUvJ0mU8vQjmLuj1gwk0x2DTTyC+VwJI0g365JKG49wBQqwN7Ni
2PLxh1oofZJRK5A5CRwg1xu4Fh8Qf2aCR0h2MXgW6Ncw5W+xiO0bh8xGIYalk+fS
g9USCq3t7fHKyrsLF994yPbyboG8u6MZpYjXBAKoL2BvotBGeSEToNifnQULIfjl
v09tyUyjvWmtnt8A7ynqAYo+0jgsULj0BgSInuEWvr/nVIp60Gv9TMOnw/mL3/CA
G7UOhvY7q4EywCkGREOy/SVIKsfbStzUCLANV9y1WUEim9FZgrfCTFfNlRohL4ex
trE4QTyErWsnlIPk41fgHj5Mys1xG/8IHtDrv5b5loHpttemXJExssZNJK9GJtvd
qak/HvlDhVtI8riwCaO7nq8WqDt9MSh7Qq8VHCeNB4PaPhnBv8O1BqsSJtI6pql6
nYYJfqGVEl6K9Wu0t2k15Snv8z+Hr8G455fDTXTTc3CRD8yL8gUKZoLe23+BCmvj
qBXx0QoS7OQcvDKB1DiDEK5XnFbG8vtRqV1jOCzKbkn90VADDiMilBLVl9HazVRq
lsD2SjsBIqWqa/82xA6YE45HrGBJRaC6o+916+hGAy//iN0jG9yFqkyGfXeKC29q
o0onCDMvwEYemhjrKexmRMqCI+p1Bu0LrDjNfjfaur1pJF4DF4e+MWYrhOg7+ssJ
0wbkpksCG6UVXWKs0GaDxR3+dVeVd/Rj5qb7u2oG2a5q/9RdUbdyb6FARJrGgNY1
GS3g3MudkE2kvyh912v2GUlQ31IGn7z8VZ1QDQ0Ghh4AcYAa5XULgj8+WHkd2uo3
0KmzHeuNup3uDhQLCM7zw1WRjwUUrvszKVlaQP+1swYEs5xk6YZo+QH9G2ERfgBR
i+Ww09BrK5R7l4GSLBvFQ5DSGfWh8FduYA1MCfG7yo9VFn2P/oRj+wT/IuWMrqg/
9Pr8d6yC3WKEhcdCAC8fQ+hoeoGMY3E4FHREnfxTDFyot7gzQk55txATFmbg2nSP
ZiNTcGIGj0dCNTpxyBHgeyV2VmfepXD+U+cEdUwhdh08+ed9eFOS8LkE1C4u2Uis
LL1Vpg4X7dZWoUpt9Fr9kTRq1VYH6aI5AbmOa19I8cW1DFNwzQ0I3HEBL8o6B6zv
rklTiwCYhjOZR6Y6glNKKbeuQt06eXD4CyDF3heEU6r60L7SzUsgXEGc0gG7TJe2
9SMnMm1euV1uPSIAkz9v0OwnbM+UzUUQu8Dwp4q6evUUcf7AiRpjLVFmfDfkBied
bcFdxqmjBN/rf14j8bc/iF76ba+WrrBz1mLqeEJonBJBtYGB82HyV1Rf9yZaXnr1
Qng61khtQa/8TibzaVWMlV0w6QspfdJ91hgqqcBPZxqpVN/H2bq/se2mgaCtXhvi
tCPXN3jhOMBW4Bzf6Kr5XtQ3zciVJkVe+5T6NH7SurIqJevuaIN4E3LqPp0J9Spp
2eiwhz8/l3dOc8Mk3kOHGk/pr+Z7tZbcOIhHZomqaA3VnFOFSwccZFIvJKYgUvad
CjgHUFWZZ4B5HJEMj1hoqqUV1fZPlMSPr2D6X7zEiWBK6rLMGwQBa9WCh/6iQkci
9qgLTTrVb6YMxDcnNUzHpvCmbRGh1YPRSZ1SVqInJRklloJO4w0dfAcgbe6Iq5kM
pVR1596w5yRso+8tNOUqd+guV4FYYA+tH7Knc/KZQ0RG3plThwOYXONHIZmVftZX
LzfwzdFVFGtY00G7znam1MHArfCH8E4pBBEw5CRcq0LlIO3XwCda0CQdL91dMAGX
df9c9Kvc5hXcA+sGCFkQ7WzWp6LC6wX+C/MO6Oqz4gAPkcjtbwZkvQhWizZsLoCY
X/NdeZJjk1zcRhRoLFWY8RtpJQAcJuapo9IVZXNdXRYNg8bB5xd+/9ZuSbmltnX8
B+eVllW+qSIY+wCuiNKd+cuEzwwOYDExKF45xpZ5mZLAKlpTyC+QdFvajDBjqESk
tul7wLYs3a1t7jpxYAaeaJeGQTxsU5HK5iMVPcQPCtYohvq7Nez+spEBQYrWsooL
30tybCC9mFmgmfS4ftcgzqbVphDwAcQhEwQ0nEjki2k7oE5fjQ06dzOaDiHSh85x
/JyOLHwxl4bZGPKaLD03eEeSlGt0P5rQ8MHeurjnH6fmWMUuLyN6+GPpGYQh5HfG
b1wYM+r2ofKguREPKmSYxOI/knwDmInfvE3s2U2bhSTfK5MKcePW1V/ZivpOITZp
BrTZjk76PvFK2oKsgegrjSNP19/kNP0EZ54S+oxtHN4xU2OWvjvfwnL3qt+3o/dx
wLZrybMa77n/TkTIdoc68I+csewLoDOzbCRutj21wcptPDWCRfUcSCJqKWNm573z
yw2OqN5GU4DQj6oSzJ9c6SBLhzH33tUIEeX0gb1GV6+XaYwh5RaMMY27kwGsqZmF
/xUu/luw9vEBXtNs8emgTcKxds7ii++xXacuvQ8cERgmOIzwMM85EJleJ3Y3gfV7
Zm866skLSFn5bPGBDwXtiy4i7+8koCnz6pQmOEQSTXW1RuBODfcI07tVsow8btIv
37kM8bEPY21Og9MHdvq32QHPFHBRXzastoc+xWNr/sOKLYxR8sUoh9nVVEaA8LZe
bmkX79yOrp97D2EN49+rKN9856SutVm1pi1OwwSDDM2zEsAjwfsJzSEQhbfJXOEo
9nNRxCRL4Xvby1UuNts3lwq2jsT4uWvAncNkayEI7O7qUfdJzlzByFUxsad+KgSk
tE/JNVW8c0RaZzw6KCxtC/Jw1u3LrzpJ5Ja7HIzJlvyX6DHCZPP97nwytf6Id2ys
qTNe43ls4PEYw5h6r8ybFdcbPekTLOEg82LhV4V7WKvQtCcX+aOiV48p9pfbLJmN
OEIE8TtAqzi8nk8lgEOgOAYvzJUVQka1ywI/SPq4QXEiZ0lNyprQY0WX/IbzeBYI
kyEmFUcD/lvJuhuBoTaaYfFsT9IWRhZ+VFHL9VoBw4GVkKH4ZPIktc2qllUOWMP5
pKxWYwle6/ic+ipnK8rjDRzIy9xdC9E+BJICR6DZ7Yamkxx/hLHDumqKxjpWHZa2
+JERpRWsvHg5uKyi/qJVcxJoMduS14/84jLYZulBoxFHv3aOmKndagCcQWYHf3cr
YMmbpNMwb9d/PW3a+NS13s5JWugdaPTJ3Y9dAg0SCoG6C4pAL1Uniu2GblwiJ+JW
d8nhbZsH5KupNd3oVpzyYbcEx0KEnJYNvJKLb5zY4T31Inv5D+OqLab4OB43Taaz
ahnjsz9PIMQZ/rI2+pXtVP0pr+lJ6UKOBucV81RbFQaqPsGmA5rjCWrdQkK2tmPa
8hvye4yuB8JI9bat2ECSVpIDxM91ydwiE3A1GUTscriORvMhC0uqcQCLssoiwpHP
desEHFfml84YraavrMKD2vmQyWT5mxwUvP8ttPytUbebYuqh9/zJvxtrG1klsokw
bE+j2z5tj/OaBcaZ6bjX965eQdqu1HfRncok8jBqFEhyWUuaOnWI0W7nS/KUjV1d
VM8ZfaDe9WwZcub24BJwsgXHmlepz8YNsFU13E0zr0ktMLq5aWRmhRtd35Qfl0nA
WCNbAkaQJxgH0aN7QALNPjPN148L3F4suykVbPGEKqDxJaeABVu6K4OGHO4DQu5l
Gx8fHYw8QwSONIMlO0ne+CLKKevr0oBGEZqP44d1MdZid1y1UZe3sDoPMDQT371f
0syAndHJ5YIPkAnGRl0rYVUPppnKtonUOq8SqgkXjTCI6CcbMIYLi8WDae6eFRJ6
lpQz0UzPPIpQSu8m3D/DY70uNAOzJQ+GOvVm90Fw2YmiezPRT+biBehulXKtcaTP
B8W4oKV/N2PazjLnJVJZegQhl/s35CcE4LTEbqs/syv/ZKA8LmTO4ZvQygzWTS6U
KfvimW8+Mp2xpVp/xVl6dvgHylLS07nRc8LxWewttAqiRSfsHv+94NDp2FMWfR9g
NYfqGtGQicx1TPo0DrgBmRhZAFVvxmMp7Cq5f6rwB3Wspupga3BiL49/3O4vWPfe
mkZr7kpB7Zk2wxct3/kPuhHli/MaL58v5M02nD4JG2r+a7MBzHjVXUePjFe7MxFC
1izl2zSXgehYCVi+9LCuoNlMtGx+qBf6bHWg5irwJyxOuiSuTGv+XqUamqCZY3MA
baIyULWVOkOFA27wvyYl+iexOInb84OVT9A2l/S788RChVJpqA/oEbxuCliTzlJe
I0ey53nndNG4vM6jNhGSBnnNGhSwxEbmRAb90vmdXrcnyPRcl9arjphnLNDab6jK
9McnICWDnC4yDGMBoFEZDaqklroP3+yAeovdqhIG/M3ko54uo4sAROyTMPSCrOta
YQPOEulKuYSfalGqQVEwU8Ap3//8VFcmcOoGFLYdz4oE4l0YrrJ68eUnkunBe3Dg
8192in515H/3tZTQiSU0ZKTbobuSALExyzdxeetN6etlH/eZcdjsItDhZdVNojxC
eV6Z8qlOjYsYmIBUzzozM2SCpO5/kTCJhZxERxrOOCHsi2fVBVqr/wvHVdB1/nf5
yXwcO2lxHT2hE2n0wIc0gXaU1Dx4V8f0Mb3057l0n+8n++sHnhPpa0Lnk46C6xxN
i8+gBm/GVX7yxZA3ppwmkgG68uj+tdz/6xTF7osuhp/wq5W251m4UE7NcGKuqmIv
63MFN4x8TZPc8DAPK+QG6k4/3WAb9fWZs2aBbps/gskNSkeOY1rq1VfjG4QZ/9aJ
Vbs8ue7Moq7vVNSkHzJz3PkYdYyo9qjeh9BiuEtC7jjIg9vIVyLb9bqo7GtZxFKj
8gbc2bCN0nROwy3ejdA5Ftji7Za3hBipvVRC+hfl91XPv1ai8p+wz2B2yaQfnYnc
SoCfu3V+TiH/Co5S49onzlTpESHyQEf6t/IKL040YzQj13naIju90rqkfYoHd+9l
xBpKGpiczRbCBc9O7/j1J9DP8WsuJfRyeWVx21ufeHWVO99t/W9vhf+yOGQ4ZZN8
LWdKCeAEfezUm/VALsQo7WJKqSbFpZ/BvvYQI4QUJ3bMhACAxIUUKU5Xowc26UTr
dN97Dnf7eoGqc42f5tjmd51K9ZetZuBjmVJI28WwhUmjEGc0svvk3OlEh6i0P0Ql
yL+kgyVU47jEx9mx8TCUETndixA5xhw/QYqQtCNsddNLT7IFOROQtFcwRptCWfS8
0c1p5mhbIaBpjYHTqDQm1uN0t1OmhwBSy0nxJbaxOFvfnqgIYKvaveOWL4ctA3aD
OAk8qmmKwTS0NHmdniNjc87GXO6EzssxQtPbMeYydfiWIh62Hr7IM0F5I+fi3LEF
BwTU8taO8ZVJegDAbWmAnoLawaJOgCnLDOAnF53oAyvH27SfYtS0iI8a8vt/9bjV
sBOTf3Dn0JKMy7CTc8yEIBCNnDUhI1cvH4JSf+BwpAEQEJ2+F1G9b51h3DVum+d9
MLVir68EcBHVKdW1AH1kbLV6aUyyO/RFlv07PihEfCFVJ9cp81sNJ/zTVq+j/E/O
JgNX6ohaddZ6oF2CNMqBlipfFR+WVWHfcEsTz+GppJFPxbyB5lhktR/zLlkMPfee
LY8FNiYblUQGUrG2jHacwdpgSJpfZfes5kM4R7cmnIThzC2rsQDkmPwg1BaWCmGK
3oHbGEVh9oX+k1ahbU2b+7jTK4HQ0iBOC5VZ5htBk+Z9vaTKyCSgM18eR7rIw7h0
IG1+pQjIJ2swPr8AbN/gpzTTeezUSpzqNbKLucY1ky25M05A7mXfZs0cbNro/vYl
V+F0M+8IVllf8oBZxmNM/yDxCXgJROFrQSeSABF0NbO54tbtb6s4NYGl65lRsKDE
XAVyfF6S3MMzIzSqMUaduq/6AeTKhxPQZ3ICfT8yIfE2A1xdxUhU/4OXoexEypgu
kSjmNgWiNrKyS4tObUci1rE55nLKMhyGpDaCzdRa3JXRzd5WZrDTbcEndIyn/Qvc
4Pig48PTEoACBN0QLTG0rWxqsOfltGACp6Rag7xl/0P19Dp8b4DycXifiYWwWw8t
gAlDpbGxq7bPmQfO1HGhbmbUSZ6QI2k1Qj6gK0x7r/cEN5xMf+sgI7TTaEUH1oDv
MTo33m2Swk/rqj/MR80x+qPlolmYmYQH2Hh1hiiA0MwDHFhVT3k9K9NzcC00/d6f
JnAKtIr1WgFo/LZVru4S8C1uPsvACRVkHf13Efaj/FFGrJ1p9PDjyeP1WzhbdcAC
ibp/N81IKWD4eRodkYenS3qYnuSkefULLjfAJoY15ygmAzcpepbo73ibCWJbrhDL
9vEaYV2x4yPs+PW1K8mIVofQS3FTw+ril8hRrkPetk4DFiJ8JfeeU1QCZ3DaFc9Y
LhkhtKVLKHHPFpKA+0WgUVhWSWWatetgNYe3KsjI+sDwgeJDb3n6VjrdmeBdCZuZ
6NGjdG/EwwDeIIiL4qjAQhZKlCNgacRLm8qaUaSiAegR+tDOApxWMIgobwLtyud3
kcEN3AYqnGBGRIHPYzlN0aiBknGZDGAHIrlUAdfM+ZSGNiGNTiWY52jC5+ClWPMr
sZ7XRWpuQ7V1el5tQYx7pEmtLh+mZbAiNUC9liXbkhUlC0hj/IXRcKyD0biQ/JlE
R0Nl9rXm6CvEPpdnK80SapPkQ1Xq7R0kEk6ttm6rF76wUX42wP8FKN18ildQ+yWR
akM7ANlPXBVO+8kjkLJMOls6L5EC4WB+ReOs+umLfAzyzTZg/iVMbKgKFolyq/mQ
PCrOwMC0ISkjesnLiX5+2h8kPwOSTlw0nuTq9ESsubUrXP7CyDic3Ky0t0mTACfT
/QDcAr6M9JH+h5bavb8Ef8pfFG0oqVHLCu+Raf8CZBb0/56WxGKlQQtlswTQSy+u
NrjtLfgNSTXLZYbNgYWgXdc8uwERmHzyGn8DD7DHtq1XErkHNdbwNzISSN9L1g3n
jQ52CMD8wRBaPSPqDkrsgG8rq51wQX0ov4nbsrRehsdGQF2EVGBmfi4IPSt0wnCZ
U3fJ3Tnsrv3vOjEq+/5Ya7Flh474hdFBhvnXVspkRLgXjwSw2mFxa4UnjZTd5Fz9
rzwfaWHu8oCpWwoyYabasrSYZlPJ7BQR4E+/K3d05Vi+z+O9NXy+lwpfS7g8Lx6o
uUHPQD+vjYiWpJJnJR6X2AB4upRisrC+2cLMMRSnnwLkx3CgeJg3H20Q3napK+kD
PirEyI1I3AgexqjG/2ZmvHucL52jFlP9sdfcy8mIoBsa0VMdu0xzkSRLvdn4wscO
xbp2bGH2jYKw7WdFMDuSZUtHSEG/jsXTzUwrvd9SD+ry9Lc6oxRrr3QlWK/cRe5e
HQ31gTAiHhcHViT0crqXZGuiebuz098NyeDQt2aqmLwR3hbNLQmFrMowgJRatjK/
nquGM+B2CHSR/eDA4CzEVgzBndozJgw32rd5N0R0567iMY5MyUOkTiw990FhwnBS
JCTeiT1wsDOR+eta0RCydVKNO/wr8SqF2wLC36zCxFT7afcTZaFhbyD6HHYu8FKd
VLpR6wAA1q4iLwviDBBXajevy36pNclIIA/zfU9PAGT3319cCdvUzXi2AqeymJx/
uxGlG3ODM3h9xFIkJ6+PW/tg2MfBPlVdMKq6Fitow4rYdAdK3HfdiJoQXBnGwfGP
FOR65oJJPpaCTXjgE2yAElAndjUyIp8ZTNslfg/HGD1PVcpRI+bEvRwnyGbc1rUC
EIm0KbGXZopznhIM0WTEkBEEXqQDe0ovjwKUBsEeTjt75wbfZLTelp2q9U0sq8pe
33M6Dt0DHfjDZcE0Cy99JETyxpoUHEvBfXbDUsPwkDchuEQXbuIpS5Rc7wXc1nmK
Wb9M8r861UADGfxq6YuEAjlTPGkizVjAOZt1VYM7CnJ8GSFB5UIaPQbTcFaDPOca
3oQZKAJgPeI51WkNiLAXn12hPt2xUBJZYHbZQCnMp9fIdGsoRicXxo7Vd05i82pK
uSN1PlfIOBSBzC/Acbk0kq995bd62xvp1X58oB6gJKJUHOfAS8CnEgCGd4Z8PG7z
D7J5ixPXZU0itk3R6pfECdKcqOHkgAmMvGBRo94O4YUPKfR6b3s3K8646qOxoN7E
LpoF3KTxCJaZ3G7JCxtLE9csynWGIZ+8SvvvqWzHKJwDWBgUrNP+IhDgFt/JSUL5
LNVXaTS+G32WNn+WcpZxRiG74gSKvlfKlAyomldy1KX6ONZLTtNeT1w4ak3QYmiV
5uqGa7AhxD/sgxqArvm88Ti8LtE/qadEHPctWYHYjuT78AHpaWf8fBGg67RJzTj2
qHm3J+styxLXnIYTQonLPXXwx0tH1a3G+lKnFbqy5fk2uOQ+lqi2Qxv2M+MuwsI3
MmnppFq92r6YB8QE2Ck9BBgNzMHuNPFhwJB4bBuesnI/tQlmDsK2uZB0hKqCjMQt
MUmPCBaDbBUWUX9KJQb0e843Vr4+zRR6HbGhaD5eNjDK7MgyiENDhEfbSkEFYSZO
9NGchBwFWRUr7WAR+43OwVjYPygCVlnyaRGvmMVO+61T2X8AGpGSJSEDmJLcV3fg
26aPS5Shy/luB1Ak9tfmmMvEdLqDe7kbwtTwhR0XY1WufwEQWfI6CajbcuQdkGOH
sIrwjyqYYiW0QDlWG/SpXtrjNjGaAN1ZkDcBftv6nisHg8Lce3D4P2hJ5hJqgx8o
Li20Po+B1ze7/0+DjSA6XhaViL2JEBBc+HFtQNEr18mlrJEAspZYbe1Igu8ts52E
lvr7XWRXcGLNEJoYJhkk1L2OM8FsoyflgcKbG1mWLUh0ScqguxH8ji+snZD0qDkS
nN5BmZS8OVzWRMXqNbDXzz+X+rcgrMl3MDmht4RoqY10A1kbVHnFi49NPm/3NYf5
2RIoEQhEnZGmLHupClJWFj0NzeLL41js5EEFRI58AI4TIjY4Be+KNnUHq0y8b28m
1t7ry1ZVZl2QjbQw1b7xctTXRXriPLvUSyP1cHln3myujiMmGZ8vrdG56rh/r978
4h4wOYsPxEeN6TwpdD2vYbeOJgABI28G47EzhvZLu+ZhbMgCXWgPMnkmMeb+6/8x
jDV8C6RMG1ihBeKNRMNPaJlcaDquHaU1DaKAFu/gOuKhLwhdW2NxeBSG6NyoHr8b
m5Jb4EXFzCvwwFQZ70GEb3GDNagG+K4gMvEB4VcSEh+rvD/UrMEwniswV7PCohvT
f4fvgFPd1/dC/GdxzHQS7zmdLF0wQkzGkLujZyKRQ9NOL7IrgWXVboYlnthlWlsO
xQciFvLo7TzIsAPN8zVG3hdb9zUyRxVB+ZcSxjI4DKkdGmgSvV6LWK28+a3KxFd2
oU+twwoVYeZyOcXr2RjUTIGNJYOS96xlBO3JGBtDwXDpOYoeGIPV9LDBtdj0WNLY
mX8+wuZ4WStWxtxNRhp7stam9zh5TUsJfWfRvZQh92kE2OM9fU41En8k0xqZJAwN
Jk1uGRzwS43peHYgJKl8xEXiAQbBE/ZTuLsvsN1hyNBsxgaDXJRIjFFxUEeicHFh
jKaKrtWl40ov6q5ddarvEQETQFcLOSFy3WcCyadpWQDZBhbC8nrJt9q55rvE3pbc
0EMQyzErrlf8rI7y1Xv1PYqyOsYLrPkZVpn52wwRZ++9oqmbosNsiQkY+lFcNvch
9xPPY4gj5NSxn2D2YgpfmlUACj8EiY0ZLvMyNwh6nOAQrNoy8NnwvRLjGLAnZ8LE
LCTR99vYUcTZfWF+I1bE6N0+hDthlCMin6Pq+qs7qs6AcVdHL6GLOnVCGi2rQPLx
hzZceK0wn9TSVIul8XJ21hCYqTa7+NQNHMdPPo/pIGfFqvgheUyiflGRBuB1VDQk
dIQaDa4dbrdjIwdyDw8Mt67un5ZSDY++GZGfjbp0ufxlyAEbF2nXQLe5G7iD2BWH
BZh/bSPBoHCgyZ3D28ZhV7Z+BbzIqdAoYraHpN5pq5fdhh7foSuw5d1q48q01ZO0
HPck9351i2m0OZ3Kwk4ApgoAdyEGz/j1Cp3ksztHug2Twu950oy45fd5Ue3+Vu2w
EKDNCchBJUXtMN2Kks1Xq5+g4UQzg5gi6Fz1Qdn4xNnwwy0Do2rHo9niRC7rZuOb
bgwJE4HrMIdpVk2FQqJKGwrc2B6oHIMS1C6UnvxR5f3QJDiMFq+N3c24yxP16P3T
NIXlp9RanWilUHegM8o5MHxGhL40zFNKwzgpIcb1nM2S4PI7F5Ke1yL/fzMktPlK
tYvkiaxa2iXHmOmGS4vc3JxXL+KS8OLD/vPND7rAtyW24glxdoWxTm4cbYtDt3Vb
HdIYmE+WxKVNWyF2OPwXsaP++WJrHrvZHc/PvNX7m62krn70u/5Xsz9/Uzg8in4d
mkFZN8ykb/rDsUncQ6EABa9ajtR8bVnd+4G9pb8NN0zYrR9Rz90mIu7tFPD9yyG3
ssiRCY0Vcbc0EGMl8/2h7hDtnK8bq7CQb9a9HrFhkb4CGr7WMC0FvxdqDbZ61e5d
WvVpgU7mjEC3juaV9tNceYbfjBUPCHsjzkz8vQOc8nl6HRe4Swv/NHqm8zy0Rpan
eMdC1uncHSkRY+hGeuTlXYGhxohWG0xJfZyXFBabzm4C+2CvePLo9xvVrvC2aC0J
gWu+iDDjGNP1gaiNhftWjqCHStT2aFiveWg7v/hrH6GzG5BrAdtEZ67cVphYduTg
MAbz4LCBt3hx9weBi7+ox2A1NmWb1pMfsQarO7rNHuXGUHfIlbAc7nPiUNn7tMN9
dbyiqykbDspIdFYweooBKmCx437kp/Q9w41qYegFKuWLPhA4LsR/JUse68URbD+H
6DZjF4X4ffeL32TNNLQ0nmySomu8uSYKIqyagkyQMXvoUcIp94aBOAn0IJaZswDJ
VIdgNiG9K+lCigdbJlywmhtYSn9DA+CjrNpMHkE8kUIfGW6vbZFRYLasE4EITwBJ
hcHe/KO6Bf87mzcz37lJXY0evlVpqIt9x5WWOkL5GjWYXUxfYWskAQRvORBJPJU1
gp/UgrzaU+MhmQ5kPxFImyzV8EQt98gpGIPfamcp+XucBfVVMurJLhvgBlQKmHp0
0UljkzIcm40cYqT9Itmlh6nZEKgbKh/ySPWXQktMu9WFVD5PiPK5AXXG/KQHSU7/
yoLXsj2uvpOhpxOgRbBtv4RpKjVW/hptSlahVqS2mTWZOTGprWoBebIF4tC1j2bf
WMSSa8VfiVYCoEZdv3lW2V09seh3leg10kRflnl4kCKTd8N3Pj2LeL9MsrHRLpI4
ZxvhmqfVAx9/IOnkF0ZgEtyPMAKhmlsGHqPFl8tEjoi1d3X02t08uTb+B12Jh94Y
W5MTdFAZLpI8u3MZZ+HZpLtSjtB7fISOYufFPxl6aDhFPiMSdz32XQB3fzST59nV
sc9oDcoCK9wU46sMbYJQ/MUbxvlRH3l7/y7dQXQBXo4Kv9Jq28hXoHO2MGGiWS5p
j9vsjoaMXv/wAY1AKCRwkDNmyDw5jxxz9sTzjpuNLmzUElpk8n0gt1JXoYkIcWPp
j8dTEWszl5YYYVSG/E+jLGGIshsDr2FZciG/0pSzpMLJWQzJddKaxemkxFlmAb2N
GwUmiYctrYjGZdNIo/qRKzunP8MOmx2q+Lopi7xVEtoJLe7rSdTa/d9AWVXnMIyj
HovFKafnmxElhouqg5VhclI/1HgYOONSqGCz82YKtYsyBTy1wwfhgXTE3CWO7STL
CxIakfR6tCA/z5oPK0mPVwpfRvMCl5fBVyuEQBgJaTSOtHPdIYe3qgEFl9MLZrsj
zoBHkZgTN/aCovMfw1ekIlkGF37hKToCz09v2SxtGFvgVsFexTrneZKe5KFaR8+d
QehXtLDf81y3iRXBn2eYpXaovLU9FYPevsTzJcopM6TzA6Otow++ud6QijYmEXaw
Vm+6uZroQyy3C3yte7OZuZYj4/2jQNYBtDh+t3WQhPwrU+Vxyas2QNPxJZpq1u9X
wH6QLFnb7A4E5su/K0NieFYTvTlJmW+jZcb2X81CTShOAfKvr/DURAsUkSPydRb1
svZzDhSddKqcLVpGdsn32Uk6aJ0KRy6Q9QLBNvUxjdtQ/QZhK0D4eVWAI932jsVP
KflnZqOghus4hFXj/khWDgjc+5F2R4tVQyPjrabPEbM94Jift1M3GgRK9P89iG2O
9IX9LgY8jCH9zaiVidWy1uVtI1Zp2RuPDJ7jmWGYylaV4QQCM1LPRrWo2sbtvn2p
VqWg6jt5wQHcdHnlVvDbOPN83djE353rylGA3dYGwBfdYgD1IhrGttIyk8End5g4
m8J51BX1JgzqcUdBM6uE9D1UyFc/j5fH2WeicF7GGUoKbjJFxbsf00ZoTdpcsjga
8rqGhWmS+jxvVG0BEHUkUGfjhTmXGrFCR8XjlcQcFyYEjgRtGSNkKDMwN7YTs8xb
qdfEctBr8OTEpDFcLk6ZofIcrur11+rm+C6/Un2vl8ZEvhuHnk92OKBBMdWr56Av
RkXCd7mHDY6JUp5BlzhX1m0lOAQaDHle8oJORkn8anEfb4BcKejg5asRB5q+BaXh
o1q75bHT3BwFfhyf4evCYstdCrulbmNIp9wXfxT/CNaEy8KCUqWHooIoZWXMMWoa
vXstCDpib/ptrLjtXmG2gu2qYFdVeGZwYOt4eNgSZp8+fLpZjtyqpM/Jh2BBdJoS
7FF0fjtwryv+wpfHB95ZZVqQ9B/rHnV1Jv/bzfKp1klKmqFpTQyEFuMFxK86b+ti
GhT+qgdDy9N8R7OQkNsWoGkbXBOdye78fo2isDmVNU5SfcdHFQpzdBW0Qoa+SALv
fwNrZIe+3GTNUTqYHHWd0TE6YbKTinltwzgT7bHdH4Hzav7Bq/MNlwbm6zBGRH90
DQWV4zdPFNaMRW7Wum9KLrHJ4YQfgtMJkxCNraZ1sxs3i6p+ZrzTDd6ZHSdKVQ6o
EBc86jCFEuMJBBR4yBS+8LvAKvxjCTEzF2Eq/a5XlAAuCErfzrK7mELTcyTcVBXH
ciT5xoeMaiRfMbvqX22Vimp/3hTt8DVTOyRNXxY2IASpe4P0A4wzFVeYUaEB7xUS
Yk4Q7pIs3F66m3O9pJ4apnhlZltaUNyDSJ3lPCJ4ZVVwOZ6GbxDDTcvWL+Nub3mG
NtrEBclFGF/kpBJcsM9wCNn1529h4939ygHbSh6JTiqYx4CDUQ2gNzJAtldxYxOS
MQ2TcVMvSCtwbs2zSXF2d2o+YReq1az3UjJoEeZcwaqYQzF7caGgS8092zuNYjpL
nXzQ1cHWNBN4LIJ31fod/QMqyiKlRbJ0sf/6ar34wTeIh+sm3bslbKy209ripgdA
TbVM9v/jiVsy0YXmGMEnMAv4b3yam65THjad68Zwqlxf/VJ9yj4P17u5qqtMHFOv
X29JrfPy0CgGolwB1kXhhDH92Q58NByJaVIFe3gETAFvWxaXay0iumy5hF3sFYKR
sVxycVN/cxaE8zpuHtYpIVXXUHsIlX7ew/AHKeFzAtaefvc2YUQNVfwDiNzGhF9V
jbbAIPJHuqnXNSMGIuavs6c/XtKacrN/renjGBvWLwhC1x/KKoLtNTqxvGNvA2Bm
EbWhWjDMUisiFqk5rM23c7sA3q8Gu2dZJJbVbU/IfkeQuBKxa6/Fz0OQvWRz/+lf
IE0DyfBucf0Bm5/gtcy2WSYK9k8H/ZNTRV8sHLRUsBYryCCL4xd2er/NI/XNVG8y
EE05X6pzl68UMkLaw/rZH6x4klgxsjklK7bvyvr7Uc/rUfIc7GD8PIkJPw75zxaF
m8UcSmtmoU/mqy0VvLsDR9TN1xSMIYUAqGtvQ+FWIkdu3Fai4wAaZMJpEVKduBeE
xwrY7ttFwM7XKBE8xKBQfov+ozK7zoZCVh3qYc389LHblTFuybYdoT2QoUf16cbl
q4VxsucU2CIjLXcWu7ImZZpXtdqf4VtOnSGU6cG5oqJdattJ0K7UpECSNzyssxqq
vNKEwHWrzXQCJCH8yUxbg3GuPR1VM8ZXo9jxTnPKb9mAINbmrHToLSLs2ojYI7Oa
HT3r7vlqWjDiWHngExFHa1yvSIncZMED/b9oklQufhUj47vhvxTHmB/DbXZFtCdo
DZF4d63ODwhlgphTCkg/df2i8z6CxjxgggBcUXRhMhwZnV7qCdzqtOEGu+0OI9CH
5FjxNPGTgXTNtCkmu2V94ty4iV2hrDAb/yUs6Mqor/8114fHa/o8HorK/jmB6mCw
EOrbx79zJYC1zZ8YsPvRSit5NgimFeqGQVn9moVgKV5wyDk12olNwDsVxbhUEnlk
FjjE2TvNtWtPAiaJvgHyyynH89JiQ6nKP2k7LQ2t4YOcTisgsfmmHaNb33N+hceY
BFKndwvErkGdGLXstd2oEA/F0AlGI4iwChmtaegznhK95RYkLeaedAFHcT3M/Mqr
D+dEHW/d6S+KY4ZOfrQHyEoWR0Pd+1iDW+5vugEa4JTxqsjgjxOuUOKYDJSsUXHT
pLnZ9KRWoF3HT9zR2le6k830Jo9ExuhE0wxioNGNWFSz/OmUJNTKzuG41614W/5X
pZjJg0aNreWDPwpKy/h9/Qw36TfhkFxv63pg7Ab3OffeBqOamcDqkWtlesD5aw3d
eKv/uN2lurpPEFMWWy+YUCKx0DAcEYQRPHR9lrPMQ2S6cIrex2tQo6+n0w28OlzQ
Ch79K1hk17dI7DfkdT9YXiAoniSVQ5HV+HxLni0lykNi5isSLk1fZWud4k4ideyc
IJEwkr0IUkGD5ySr0G1hIg1l46r6Eu1oNMjx+7D3IgTJhjO3m6LiNxAQ8kVHeMrL
s7XjIXYEXbUaTPtravhWRcoH4DB8BDMw/HqSM62nZW3+Ll4QDwJa8YTN3smM4ggs
xkUprmGK+wAemTM+VhncrgA5evTYZ/c3UOdsQIhSNn75DiKRVeQKp7gBEDXrsDPu
PWj/9SBzQ6lcxuFQoe/Rh2uC9JO3BJl8gNB5VOpeAuiwKyGXRzyguUe3eoLRXO8G
BQZJBzmFF7Wnh3XnyiV+S3WMQbyAS/iRW23Bot3c/JVUxfvzmd4uoXpPTptT1brC
9yQZq/OqPJsFWdtZv4g24DXKnuqmKPubQTOGLNZhzUO0su5YCI/g560yewpSgzkv
xIUHfcX1rPl+IX8izp/YCT6AfCzFYrUEG2lyYZ2zB+6GygY5xPk+WJ6rfIXNAa/q
V91+KmOJJn70pVYROp5q8hGlv/Y3U8dAZttunTAIuQSJWw+sNHUPuif5pBLEZ46w
cz/NtzhHtQjH0iWva77ciNAyP+B1n9JfZmk6DRf++1HR5cNEjzOvrj7V25z8gPVZ
tjS/icpz8E4zmF7Lr3ut9UPsY488iCijgm3+4NGqf2iDOnlVquV/DWa5B5bfB12o
HjeaWrGFpujt1+NatEVcOfPENXJg2KpEDPgC45mnlgiyU4zBy0OKAKYmwVqfiddQ
6P+yJPQI7X1l0lURCFU/VoOuXgxj8z59fc0ItqTiq1vW0hrWtE49VDPP+t7tw8BR
C8WJFnGXebc0G5BWDHJftRH+vqqGY64xVc3yFpGbORynr/kfHOOAQIQsVs2nusUN
GAGIOm6D4QHbPd06ESQsNXvHDjredU3e4o5DC/2QbNnnTjKymPW5q4rCxGVzAy6L
MFXfKzMs7pQgkHA92oqBhF1eZWhhj+z3MQCYQylbVTMP3V+9Qj4ZhfaXVbHw193t
go8Ppg+HwnO/mIpjFCzKed48QDib8cMtZHHUeyAMpumoY34PXxD8fdqPJv01obEv
TL0W8RiVp2o1hPFs2t+wfnE6PMa3iaI6hL1+LdHuJuJTxPN+EOClx4ECX8L8Vpsl
FcUwmOhs8aZ3XxgrzfM4Ysb1W8nsSYWqrf/wCCkxYjRLdwa0q8NjGKfemgXiQDm8
GZ70GPI1tMyugFgq+eBf5KCc48juAem2Im2Nge84d1RhdhPMB0BnifLaFp9Mi5ph
yTIv5EkKHo63bu+F7Ao+jnowt0P1nNPB9IDjF48PSZJbsJbQVVqZ8fJxnLRvrpOK
kZLXzkwJUHY5lo27wevPGmBodYm2UntSLSP2ovqyAYdhcsXdob65U3kVSQ044fxa
V4ZLAu9j4o+R7kwAnwUDSAcU2JtiQAn5PbsU6yU5dRWXCVatgHdx1lJxTM1WMFV4
gziduHPCvCP/ohrbLAH2xpF/lgU41j6suR1Wg4Sk5Q/l/hMWgpZp8eTdor8Y06jx
WNQePLKkEzUFmsja69Bz/SKKnyvnoaU7k4YTznXH40FMO3kG+vMOYHCXOqulON5u
MNUDReOP3OTzdot1FDQxvPOjj6XRmpXVkZm/+sM2HCfWUSF6fAeucH2YmlesUldh
8XgKB7nWz71DcmcPSJ8T+pfy4nrGN6OcIObQ2CvcpO/I23JON3MQqNkjTYIPwXYj
NDiaZLGjAkV/QQpCt0m6yxKY1d28v73DIJB0HEB6WVq77k56CWxHOhdyzrsMMiz/
NWEM5dnSGa93n8rNXoSNUlmHTPlSQyE5C+2BEocMDGHiWXkVnkPixt5r5e6WLVrV
253gW63qTJfFXpgoTk3yhE2xE7bDGeKqSG/UOz8ff85/wxY0Kl6D8yoB0nra5G+9
Vee2e1tHHPAbblVroUmihhXDdx9Szx/1RcHPP753ctQNPsNZhgtU3uST5ES3E0si
mzpYQrOI3cA2+1EuUxYDgrBKFi+U/1OY2RdFi1TsVvtJMRMrdwq7jh+lGKqq7ici
QcV2B3Nbi+l/YDAOuL4LkyS4b2ytSq2DsEO2ER9QgfLwsL/rGuIBh+ZCn4QoOdVN
V8E0EwmPED7rtSTJbG5qlHo/p2jxKYicFaK7hmKgJOCGdtlZl/Ii8P2nmmZ7ooj4
zl9hg5NqNp+63qDvvDSEq1F5FnIIBNWR7m5ixzJJrLtCf3YPrFSwWmbvPxyGmk1D
mY5iMZtnLK0ztA9K4++7AvNkkFfGj8rShHtJ2nlrrlvKQVUrzgGPK1alDv2nwCKm
E+K/A7Zfy0mOgDq9Duu9OJpip52dcf+Nz56ZRmiYGHUF39xUeXOpoFZAqYhLBtDh
uSmk9V81CIXMG4/k5SbZxVwo2YO+yLPnLOnFeQ+iVATPvk8z58igDSOnUFOv8usB
NiNr3CnvCev2JLT2GVOEq77sacEe0VKUnokFTlfzTSKXCvk7YMRaO6oSp9GCif6O
QaZnjikN7Lp5U99jSS3wnBfpUOMcxyFXR07lWtV0XSNICaSoSxdUC1qyhYgSoMNe
xqGZsj9RKFxFMw3ILNLUVR19TXt22ETsOmiV7tJRTuOW6Uo/g8XYGJh3MDKmAaYx
UC70tkYg+P/fDQjLYX/wn24V2JC6RB4Wz2olYh8qywVWqGaKOX27LqMyixb+6NRN
BwSm1Q9bxxXfIiYC/wugXlSC6fTB+MofSDgySFWV3sGUf5Jc2efSdcNd24mN/3m1
U/+OvZmcox4QCNMNpkOWESq3u0HBLWKdtIilDLdXbu9AUw02cd5XrMuvKUN5V9kZ
pZYSeadW8TYUAeSgPJAeSAd69NIrVs205HuxenjwPI/9kp2XPqaiXU9jAQ5rz+QK
/otBPc1hqH4Q2U/ZnibxU30Kk86Y36Oo6sZ2kPtcRs3lgOM31y2bS4vTvUGawJcK
q3/8wF9ZD7oqZjrjNNK8B3nAWQhjX0fWfmmxTtpKGEmrOC7orpXoLrSsI8PLmXEn
WFZeRyOIVmGzE9x4stP23/ZvBGSasqASvJZhQa10rePGMyP4IHjgQU/O6MGKWaOa
fz3/TJuNM2ZQsQs+e5SivVZLi4ZKuJfIs+5qABRvVX8aO0TUdhmjVXa623I7JdIf
R05ozKx/a5qxNyUQcaIg+LwVc7kYBYlUez+74sOgeJCqHwTU/mgsDCcE2UpN8gDR
sgGQ8ECCJl7RE21G5C4ptHOu4lQjkfJANihVTP1zLwYpRPScoR4hNsi7Ajg3FOt9
7t8Z1xjtPtQwzLgr1oiwAzkJibg1uQ8cc7i68ctRs8MqngW3CBMAJPWUaciu8ZPx
b0fsp9/KgNWJHeTIo8Vy+2mt4dCN7GHd0DDoKJm2CK3Fkq2fUKpUaS8uDdyU9Hw+
Q64JDeqnGzqDhM2k1dD5wes8AHKSp86Cf12aRd3AfuBSyiOxSpBOM/9KZjqR48rw
1l7ucQDsE4RbAO53WxyjxzEwNlAOghw1hY/Wgh3uRjax8PhOyQXdatKmABRjqcek
pre0D6/t8BDyRZPjXU3qaAjoYYUghMiTjpYFEXsW9I88gZ8bvxFrdaj/J4YfecfC
/UebmFQ1duEU+OOYmcARlN1yqAYyRPrD2RdgY7jzpYTT+UkKZbrZ5JtOKExynTgE
yiqX/OKHzoHsBkEyZxdwvhKasprsf20DRRzEkB6cr8xJsmQZ8xkK3RkXfGOt0lU4
X5ss+3iBqUVQPsBkBg3A/3E72VPtUPHOGrxScJbdxKZA3vehxj4m6ZWAenMixzo/
yVxWQ/IfVG6lD/U10Gf/jb5zwcH47SVKnCbLP4LsJybNb98oxyBQ2RnDvCDC/VpZ
6XWiwBoM7eBZKiEOwnnhxWzLh/20Df+rwY2LAxPecSE2keOqx2o61ECmvRZx6N4F
ZXEXWmo9cm/LCRWSo3oRYSD+iWSTgMAWyPYkv82NDsHC7Y3MQDcjkDpSVgHhn6Tt
u9eZybA3D47ywg7HM1UsuGptRqngQuVguEitAqTORsWbXXdHlBfTU+ds8jfjWD0n
bcZexiD/mJqfFTxhllt0qe+dLih2wxtlzCbh+BuxLeIKlhURDpZB6e8EKQwi0wmm
n/aD3QvX/syQXTtlMrQLREYBejURr2BcEhi43PUAXnCluhK9ye4NSxoEWT5Z/gpH
REk2kVO9llim8vMW3QCowguqgcnRRknCsv6D7iWqdyaUmBt9MVZ5xqcbVvHdl7u1
LTHpCpcZSCZhxLWeHsA1zfoqWgCxX3B5PG7PCfrYRZ3OFKTlJSdefBuIudNv0FjW
ppmsLQ30gMxXo4L6GInIeEEzDNji3W0B2i5hZ/VyxV6zYsRIXnqsq+1TXdpvFTdD
1+aqRWHk7OdGK6S37hDoBpHVMDWkygQDhwXpIeyyCF6td6wwzKMA9DKouHhOzEcg
6Uf+ga2Fsy7sGanP++Hf/eVflUvLj5V4SGRLesH2wOHVNxwOrL0H4394/GPdlXb4
z+5Bml2/VvEeqQOSLwqqZe9MqFzizI1/gEUOvNw7wDOHUZopjQdW/xesVVwH6PKN
6tsw+Yim/aQ8it9tydJdugcxoq6J2Yc2SZ3TBGfGCXq2PjFN8e8fylfGDOdoZTeW
R2QtFToFx63I6wB+hKwhMkY45nWKSdG+iDhSsXfexCbji/J3p3Wj/jNSY92LRqzM
By0vE0Z9LWoSRTMoB3fED+VTgYSEy+ewel4PPlFDSaJICZe3kbTrQ5jyDjPSQtH1
jK/kmBmuLVkiD0JVb0SdPZVkChzh3qu3Ftnujx/1qbyx5qBm+ywHTvvYxRFfNbDG
d7e9RLktUOaZVdnlZ2NDnaRT6UMfwxf9IjaRfEwABv78sa+gTb+dJg7QSOZipUQo
VTfBQoX0049B03wyhx0AR5ZWuqLUrcGgSK1CCR/udnUMQK4j/j7AHH1xRh+nt/EM
9ln8wdkZiWsHByZKqcto9vzZCVz2lgHMkdrl/9zs3FqMKB8fplnmi08JgpcFoLsj
t0EbLTVKCf46XzkSiZLUIb1vW9lexKLf9o+DdO9TS6y4yN72OIARGg/D6TpeNC6q
rZZe//6Hx2Nhi/FseM553oz99LVEBQ7DG5OrnRWsd8CQ61sEn/xI5nIDgSFRMdL0
K6TJ7/PmyU/3Y/Bx6Os7blvFEGlzol9shjlygwVstFzBOkvzMxHqCvhxlC6oJ6R5
ICi+N+2G+x7ViR5qa5/yDBsGVCYVNUGJLCGBUKFfpUZJJiKqFIMcQDncokFUhiFW
87ukaJdYoZEKBpatHo8tQAxuJR+/LvSzsBMe17iiXCeIWS2YvppOYl09q+yzGDPK
y6M2NlDHz6ZMdsNwcmGkhKDvSZF0e9Plwdj3+R3YVBVZurYLP9AbXrwtby1M64UI
17vBdhvpeB524Nb/ePDUb2qi53n0jl9uj/mzwxVBLmaakoPuLmKto9JGSitKwDok
pZHyJwrKznd9UQAv2qBRD6YojrfEplEuw9aza/Mcsc8ZRVXp5WSVqVkAsRtrZS8q
xtWL5Vg2fFA5WzmYf1IMZs5AgNzRwjGiT2Bs6Akkgwdgg2v2Wk81dQRr3519rhrx
MCTXz1OXIczc6NpFG7u9R9IhJ6PL7Kuaj+xH5ZJemFxLYSbTNx0euEd4cqHhTcGm
rBNy5O6uxfT0uLhtq+qND1VTufzaCCOInmlLnCB3hqggKWdOPLSi3150/vnA3140
WnKDgc2APG08I2xE+afnH43Tn6ijlHVXpX9XZMIwlM30EhTP4rqxSG9yjQUorER6
XV6/GZDqUOS9SMfgk2+QgK72Grpmy9MvjOmH6w9TZ45dHQe5B1vl4H+/Zw6dSiCI
ZB4F1/0Lmf47j2LbH/lA+wFFr27hJrd5hTkk7fixmosnoKgwmR+AnabJNlNVT2S/
MqyRP0SMiQhMhv2iay1DUUV5ldv5uyLt3DYLWYtxIxXZfRC/Q0lRqhahB/Po5R9E
sDHFh6xgdmL/bKs0jSGxj1gG/LShNhLhyeUAVFZGjDc+LFK+QmrNXTZRxKoeTc+4
f6h8jNpp0ExcOMPqS+qaL6/be85C6D71JB49LMj9BPOpgwLPD4mid2ikLTuR/2aM
2KWMCzo4vT06+5bTbSM0PCIbDY7OpK+3rQALXlfpfHfyg5Kgqq8xSciFLEiP9Xro
fz/hRxg4BJpki+r+Ze5djkq3LRjYjRJStuk7XJqyuzVYsoJvOP5Go9G+zUw3dS6Y
8INgntcId1VgzA00OaPBEKk7u5lHapf7qWhnawOWG4a0FPHNC25WnEKgo3doMqRO
aBXINR9ITW6kOZLw9NUzs/HGX6VHx97fB1k3t2/FQ4s2guN6k7Y4Arub8nngVVIA
Z0E7jyLMjpODPRkzwnW+KM4arzQPFRyKS1jnbGNa5BO/0drDzTWhuNIgHbqJvcid
R3rT5xRIcEpSXKyPYr1u21f17bN2AqO/8CHK6VM5wbUknDTSHHjiB1DhDWuscjpj
+J30sF4kUceRpWKc4qNTGIWo3cWWs5TTXJz0XaqGwjZ7HHAJbVIvrTB+CBqxdt8v
XLdyq5lHeiJjRXqu1NCPgDQy0ITpmhFuLurjwL90kf+Uz26xNjvjYHus8+GcWjy7
0kqEqx+/jnu4BvP//tqTnxvDl9FtetOoH495XmsMFdXzemFjejxg1sjG8YDj60Br
w4hnUxLDV+Z0s2T9ZHx+EwVWrX4MDBTzZUEIdEWXcHtdGGf/Pau1LswdVXli435E
TboA9wVaGTQsTkusKIotadi1I0EvV9+Bm0hvYCDA1k7x8MiWgBg+Vqc74Js23A+8
OUoPDo5f3yhaVJMbHyJ8t+6Y6OsykCFJdcwoAGAlE9zs6Y3FqqjPs3YgZVbbDbFe
qBK2XooWRtgL6ZsZe/7AnoGTo6I7BkICj0StNx02IyPieM7LFLKBuqeHeGQLIJ65
iaktpgXRMD3Wxy/gjJQf5Fn80P+zeURTTrAFQWBUGbDySWfBACyVHwzNp0woQlNG
o4TjozooMUPYawuTFzF+GDmzefkJ388TV1la/6FFD4D4PGFmj5hIAAYy3Vxpxy+P
p+7wuSxoaZW0YO69V+EAvH7OKZT9LT8LzP1SNcO5+j/rkUn9No2BFzWsjqEezwTZ
CRBmRqGVqCJKk1uy32XJQJpISd15+6Iair3Qsj8tAZ0m2BBOUIEm1LbeyIq4mCRS
QouBzffl1r0dVlJXmblS6qXHCwSmVNgB76KAYmFhL0MOy4zKi7gyXhqblVICRP6K
rGZosVPy6ZKCAcMeq9BDXeZ5vNspcDU0RKqjDY3rcvfiw68LWVxoCEpOfZBppUp4
igJ5/lYioh/nTZB3B1Yaqy3ZFzKz5KoKy8XGdKaJ5AsqTn8G0KPIZSI/Hs8QFroi
niZVdicc3ulaiQmhWMQq8V36lF8HDB/GzfqM/aI4pT1uYpr1l/pBT/ONZz4wpfKY
KU7Z5pWaH3HGNSlYkmjSV4Jhxfgj5gXl7wTmHDU7XSlw1dXoMBbfQCJlQGHKNnib
LHMNO2T1BrhGVh6IK55b6H38vl6lWYDvJEjJ3cte0+8FT+1M9uodolFGFxpQ/vQr
qGkhyaRA+WK6IEo2ZGPFqkW0/DxTeUK+nAB6CeIvtSmFckBjXEJBNGOgcWbY3a7o
USJ9bUl2ZF/NvWKYPNwc01jAkFrNnlF+9HmmZHQ+YgQAGCW/bAHHiqDh/7K3B8sY
mVZxcwV+75yqyRRNbM9Qqtesm7o0SXTFijxfiQWfTPlloXNaL8HOpUkY2uQd6LbR
sC5+bYuciYAQvxcGhlNMEMy04DLTTiAbcoRG/LRbazGWAuPXrapz8bHM14SB/nj6
6qjexurst3gvUA0KGF8Dd6LY0/d1yprKfuBCeX7fBqp8Erf2bgrcGr32sAhVidSc
vXpK5x1AFyaRqE+o+jG0X6tE+473fCkWZPMos3j4JQ8UlxEC1e2Mw9X6136LFEv3
hOGJS+sqPLWsz2UZ5cm2Ch3Fx/iYd0qC83VAdniuPoSfvENVyUvVuYji9xnkRcb2
/b8n8HmnbdcIB9VPCmDJgG1RSx1km8vybPer3JwQl3A721uQIrL+mhvWbSCsnEjx
rll4HcTMS6B2irjfEJV1mq62wMNzZjRY8qGIiVBVEYLF/lVtbLQZ6/ICi4DHLZRF
3SoVRT7pK8dbiNr/G8hyDh/ZR8CRYEXDn0HN++FKBZBpC1bNjk3B+s8OnPMkUJ8v
0S7tG8k2Q+Sn2qQhnoRlw9LKKZgPnvEBrXZ0e/obRth++OuDb3ne394rFBCMzOIJ
aTpiFaijrIN+3j0TcQHxrHAl8npIfx30hPsclEORFH1YXDcqqEvqGqh8mLw90Ji8
xe1l0iDzYE5KvYM/urtPYPRf3X0hZhpHjugbIqRQZAbCJOy1EeQ0coHa0fm9rC+J
QxIi5z3fKugdaYMGwJ5Clcd8kD9SKc0NenWbOg2Y4LHl99aSf39/L879M+D0BLCl
FC/Df3LTA6Mv/hqdJxkdXjUyCFXnElK8S4MEvJz66kSVQ6eyASgG6+L4Lak4KKlW
m7Rfb7oGjGqnukXGj6IWirMwsJEsUXnVnhyGfIq1na6DpInfe6j0IxCvhrIrF0hm
GrScVJGqseBDesbyCgX2XHJC+KrLO/J3OFqX1dKuenv1zyFYfF+jEgue26ampH0N
OPpExfhPLqxwqSBEGqe6h6RkzrXATKAvLjwCBgpQU38BRZmiophZmgMgaiRCVqTj
RKagay8sWLzlpHMOKvui3iUEz9kEADP1qGvg6jZqa/CnEqimzKuZ8ic7pjfAzu1x
fGrs2n+qenxrfvDRgxJcMGygpDaPogBlhcYH122fs/J6H4zgcwgQ9wMpxdjdDPv1
xt4Er/J2qg4DWYdi+5psvbEygf778mg6m5gvqiz5fUSZyLS70x5dEaPBsJJktCmR
5TZScSopm9cJkQiHS+Z2jB0Dxy4acJIbJt6UHSE1nuom1+3zQlRnEz5TYy/uB7RL
k7W26rwxLeWQGoldL2ip4xpZgK/qKc5Dq3tRLN7xBF9PHQ3GHUZU/3dcbbwmHuSr
0bh1kNELNXfjXL5DD5khVNt9s3HUfAE7e30ApW8+keC4qzbwarpMaJYxb6/4vKaO
v3yksYUOiY/ZaQaJGbomF+jRpwsDQtO40h54owriavLaMTu8sLfwVXZ4PLmakOLb
IMR226wlVnSiaqxUr+qXNrXdOZCOXJcPYqW4ihiHVYSky/bSCtXm8Pax6icbbDTF
JXLyzkycDSZ4+m9RKFiUcetLcaRLuCR2Iz5f1ldcA2fzmT1Rav3D4zPVHad6ru56
R5X+fLUFLj+jH08HDXrCNaFLZKU3Zm7KeaHGX758XEDsS7unU8KwPV+7Zgg5PMGd
SU/OmbaP7/geTtkLYzOo2ZJI39HqZw3YQLw6e+yU5/lo/ipwgpfTmh4nZAOHDi+X
CSMKQPCD2RM2IRHsXJDbZmZadCVV1K4vakceaV+YCymF45wHai25WRXSG0o/H53y
GDBUVRmXsI+JUvQry1KIw7LfkQ9IUHfrP+7g4um87x45WEbhKRm6cx09Y56WbR74
vfdDD3PrEib+oNEg7JnfBBVVR7CjNGVOa5UpgbH37QmqbsV8DbGnA51ac3XYBQHD
nlQIswD1OeEasf5wePmGTvMBDH8pKJbGLVew8RLnxzeQ36J2xQ5bEErQ2rJXj8TR
7U9eSMpez9PI9Tq9bLudhS6OF72Ckx1emhv2YTRIgV71QKnIT+WUEWtGfQCu+OP+
GZDZbE44RUWzhPnJaDzGPwHMRCY/1wQiVSApAOCXMJWpeME5reMs3F8MTaBycbew
FcEZ/Na3ZvVmlvEvZWZqT5Yvqk2w8O+mgX820hTgmDNwez69ScLLxIcNyCOn2FCe
ux6olr3bGnuxmpXD081k60fxAgIQ/DsN2MsTGWPpMO7uJOz4hFZVBhcxm4YK2aLm
lBuat5h2dv8sW/R65eKsI2Me8P0GfzpkLMRa5WmKJ3OgUixKdrSnr9cJFSmM4n3U
E6VUW1PIvDKAFhSweT2wDr1IlqUlGwEjUBnzvQ2bX3iVVzBjUNeVu4f/GtfBJcre
X8Ii0QnWO9g9gEU74hqi3w+wN0p+1pFrkTkt9ibHqiAiDc+fVcVHJ+6tSa8yb+NC
vgsoAVlClZKp4FRo9C0FWSwxZtgCxMv5R5/DxMH2KJwXn55dVIlv2gjcOuK8wIU1
nLc6Lp3N5kPV6QJ1PBXYB23jCyTRcEYwcq8biHrsQIgIUL+xGxxoaO4JolqeoCDU
xwkQSvgbrLlCnS4W2+Tb/UT48dAN+vaoIJ4caWFRJ3NYkORMwqAxo2qJYazt+Lnr
dm0zG78OWR6SoTH++AXJ9jLx6mZHkg58Q2pzrJLDRV0IDSXIMorYmSuHXPQjWdGK
j7N6op/unf7vp1hr+qczFpuKxcH4Ne7Yu1mIlNocXc0lk7W8mKcPICxp2bCigvZr
j4gotsjm9sKPIGs2uPReNPas2Jwp54U0I0Xc7monILQZQJaNPkql7sRIi3vyK6OH
FOo5nLVLyIL2KSF+aHoebWE5AUYQGjtcHyruReb6/kO8juUzkKAw/fPLAP+1Zho9
Z7swhVF37l5OaCu960W7Gu7nVLmFdF8zjXbqIn71G3EzD7kZpaRLn4emBEJPuVVU
eyKQvafXFWwhAxGqoj/mgOQaNXb9JZda/ckU/JS4pe1qM2Kp0aoNdHXOui368oRI
tFmVrsmJzlvqHqwQbYMX8cox4GTjcNlndfwelkahoFXnRuOTuvPocpV3NUd9vDgw
toe1e4sfqnVlbV1H7+jxJfyrwa5SUvuua3LJIjgIUl1tww6M4oqnYn7G6k/RVdUG
mHWVDNweG3q1REh8nPNNJ1+qhL9nInv2zjF2RMuk66uMeqxx1NKZG0BkAeHOvCrr
i5WsiDbJ/xW1mW3EssggYsECcw15bRCxVAdnzs95RE7sXtftYkgqmHCNsebSpte7
hAzclvon+eaHMUaiT3tXheZ4m9ridfzQKMvBFsscokes4Nj5wzL4S7ol3hBZand4
su3/z5XwcyMbq2oLsTJ7yp2yzEuO0sCXiuTb4NUuyY5ZedsUp4uRsAKNbT0PWEUS
H7PLAXzlRkrntFewH8kYmkIY74IpIMu+HX6pzY7OA3vFDsxeCmf8ScCWff295xAA
A3d/4B/C1jrA9WfkrLGOmc9IPEA9/uJmhtdb6umu2crjwe2xWKFh5jDmcAV/NY0S
4DbaiWvCoz3z0yg4mZHDIPbIPNsM6Fn6VkUfyLSKOXBIYE4Aw4W5yPeu1wMiPCcb
nmTx7j+9+2P/YgRXQ+v8VRbecv8GHYp+BB8u5BcYByn/rCZmc7a8drZnxlFaW+PR
+vsJ/achwU7Hxi0g88c8uLpGa7Yehchlt25k+n5rolhOm9rcSZYEJqa0x4ZtOeNH
Zs55jRY3oBeO9SJr4k15L4yTjOOM7PffbaLQsw/Fb3sXdfrnsFX3UQinyVgZMfKD
9NM99rqqso/k9BoZo9dcbJI5wa++OMpbe7AHYyxXnqcvk/EicFvOLZThVyNxrlA5
KTprIktZFx5Ehwo/rXVWgZM6pIW9KQAXhVSsR8zhRyQfhGYdRZlE/KebWhTnfygb
dzGpFcFStnG5yRBNxgvqr1CG9KbUZPG7uzbK8Llj2vs5iHKHRDmkJrECkAL5tCHN
teYjOFIH3PYk9YZjL3t2MPK0TarT4Jzr41BnanLPyw+i/SLRV105H0yyygrbD4tP
O3mh1XgIYUz1/YCYUJsrKOvUj0Mw50uo0+F5NqRCUsK3PNgSlqixN7ANa0kbh6aP
Cd1m2SeNNqDBOYC85fxckejM0nbPr/jzb8qnIuQHuw/8/5OPsNmXkRFRbLDqDcok
1osAxs1neOAsdL6MHtpjymNlIC0EVSnTEH/AyeYqVqW0ZER+eCO8Dj41zcyKUGFd
3b70OPyr6bhyE5rDLtuS2Xg8vLerhu3WKlxqSVIuheAUygSQETLaMPAA8MML4uSS
/yLqNwXMAWfrYUuuCoDV81iRmcmiZfZBf2VU7nBh3qLjfz1lRBJJULi5/cJtsS2T
C8FLYkot0NFAzTx2QI584TY61GcbUpq3L1KHfPKxt87Wl52IJB/+PcMIZFg9Scbl
99fr1/5OFH//gU66o+UpGcrk8WtmwSp3soSM74oVQS8Fas2mpQfb+WL171Rtkbx6
KhL56apq0aynFyBFl4PkkoSJwaSIuQyH/DUHCr6hismsmSuCPJMG28/x3D3DNnIU
IDtm2GLfZTGpReOedydj6gog8RZtOUcSmJyqx/6xj+1ykvXA1dndf9RDmo9Q1GgG
Hj88QtJo0OHC61XYkZGt8ts83IwqKuBSdbmAwMEjjYcPc096hHmZYVzUkuBJak8H
ku+R2ovxFVgHD2RsAfjWXrUqLCJQ0HFmYhCs/qtzpUwXrho6T6jsCgQ7BsrUL/gz
g4xjiT2+eBQ5CudRTYSUV2hK7FpqFZG9Sw6rqQweJyR2joR0AldcGf9QY2GuQnxt
V8gVR2xJMxTjKh1EyYWvDurn2L5rSBsMhT7uSIHkxkq3bZPo7riouqAOBdQ59sSq
rESpVNcg9gcnI0BaMVTHtilBeUPJBDX/K/zM8vm1+zaIXq+BUkVIMtXmLwKsNsx4
2RYEnhydfEBodmDD7X5Wh2iFc7XRAGXBSysdzD66gb1JFcp03xJLdx27f7LvM3xe
zeiP4e5gSP3Me4aYff9v+vCugk/vQM2DNWlCeUDPgF8tcZmOC3r7/dbEFH9K20PN
g1kQlaZZSE03i4ZxZk43GCtxz5aTTdFF8jnksrzSPCe21lZk33RMUnylGrACgPBr
9CsAUKpIwgoCheDw9mblKjzB2u0h0nlWVmEB8gxPiBi9DnZV67dQhTYo3ARNSYA3
+hKJj4ZDyTEZzgCCnhM6EzcQ2IgAwf/WPlQEL3Two0vwSA4nfzLWa89e5ulw/tx9
QHhmhlpMixQBi6akdu5FkTbQ5+NJiKBLvSTnMzKKqnMUyYfPFoCisO9rFhZ/FIm2
PvD0P638SVqtCaTmin+yhRC9OgYlUprYLdyodiZ3aeQwpqKk127lQQScGMuZJclq
ob9uB5E2AXiJ9354Y7TvnxkI7nAne1Qs8aoVHH762DhNgsEUhwdJ8fcOZpl404jn
MTYQrbkxTd5dFeOhsLWcQtZ0jfzivS5yT5NmnhAsnnY6tkssEMGGCgfYnqlYD2F0
i1IjRf84mPyHBKFBz7Vx00p7XezWRli3f/ZTl7ogBaolDuZ/Go4Cvt/3/UDlokik
QmkiQe/Rpgnmqa6OztDVGGstc525l+pQn3aj0wRIP4foO/k9P7x1xatsYBRL1gyX
JnpiM5h1KXh/FdVhH9w3JSGfnCjIk0YvT8hTCZYCzKZJDOoU2Yypwp/nYSANil4b
aT5u4lBmS1WMgdWZNWDHfExuZoVTgRMGX4jMLiN4LA1oFX9iEPLHjMw2i8bKNySa
zmnzP5l9CQ5OLzUo5PnJcnzHtdwW7VCdFCtGOVgR9hxBkO2/73OalnNZuG9dCtV+
9IyXS8I030qRLyVHnmk5q5eu8QLQJEy9twx8q+rSCc7Fgc0Ut7FGExahYeK4M8hg
uL5BmzCncsio3lCtp2LNpCyRHoy38gA+Pv8DJfhn033qEoNpAMmQ2EHzN8j3NA+F
SmR2317xMIFW9lQIgNTkfuCIT2Dd1wmTzTrsPdc77qrcgCLqF1qyzPPml6fsd8o0
xpANirn9NpE5iyM8u+tku+ZQkXYZZKE+VNGVO0dFySIDFUa7I8DdkEuVmhrPCMjo
q9YgNacU92NZcgqjH4yXDs4xrBChoeDAj3UOF7z6Qj4EMtjwVmDAz+52Dp7qRPeu
G7v7e+MjFzVM5zhZCAoOzAHSfIcnRa0XFBAMT1zZne5fyZDjfGgo8MB7uB9hNUIy
6Qo3TXE+gwBcPYZq+RBForAMmM2YFUUud4ne/j7iL9er3TqeauFb4NupHbaGTF9W
UQH8IreTwHxIXwCMya/trqql615IqjMyeqXTxKK2/MYhTYUVY4L/cHtMtITbRRKM
ycLV3E515dEUKNv9CvT/pcVDrtYPc4linNAVTNg3LlZJj1PiQbIgd6gHalYdxOfG
yoNpeMsmwYFBw0x5VfXuu8GsQ/luKghYg1kbSgjQflzrDzYvcZfCz4wiafAYjBIi
bViur3nDfNGbL98iQWDKc4hwG6I+eUmPruRhIaV2bVVqfVhuie0S1tZffuBIEs1K
PH21w4fYNVGxuS349Bgp9zpH58RZNs+JsUGZ2/4dzzI+iOaaQJzBGLXOS4ydEgLS
bUd588M7Mc3gyMmT0KDiyWt5bGOKTidJM4nfGWgWTqCZwbqg9sR5xHa4f25IAVoR
orzHqmn8kc7vJXgA9NIxD2tASfMOdtBishZxW8DicPXaB8NS2pnhOfBNiM45CzBe
FMytbm/Mb/qOWcaoZ1YHmUlKxIZ4bgABLBnbOtzRkh0V/YV/DDbBjpdNOYj0pykq
hZ9+6vcax2dB0HlRN64sLVKEU3is9LCYXyJqngutpEortQWWYnRBbzzgI/e18Onu
AJ1XhdCQ4+hLHjSS5qBBz0a4TONDtIQ7ZgnzrJx3BXt0e+ts1BurK85B08lRShSv
jQKdKOpE6odI8YZm8nw87PYLRDKkzBIxCKwF8yXPro0PrvVQZJFWxKi9WOC41eZq
uBkg0atHcZQHsUadUBzksLhDo4QHcqW4zYaMF2n1wu4SOZl3kCMZ4X5iCMB/T6Xu
8egyEkOuUvxcJETBLAV8iPlOKui9gXa6Az1ajGhzWIHl7uuf7clD1N4jCALFd4nR
SuGKossNPEqhOSs08RnE1tdQTL080DnD/AGzfn6TbVTbC1P7B4FCzrFhvgu59IG0
tWP03fZcHHC+RtI9mELM8sDBrWnbvQSgS04+P3ikwjmjWyIHOWCS6Ko/MMR/j7bq
737Z7kCabOO2W+sIRW5llqJuzAQepYf+35k407ixmE0ZH0LQ4aCjQs9QV3Xarz5q
MadogCJnNWBV7zcuCgEaDdTsWD7XswuuMDGH3bb1tHdtI1OZwaT6LFBKekAbtqds
lNfZfZAWbOAfl2WxHb/vVGILOkrmZo+J+OYLIlVmjnGe6ZgEhRTIwzjA0oK/+31v
1jFiHND1eZZ4JWSiWgljaRbCInb4n5NfP5TtUTuHyg9jqVerIf4gtauvFHH0yBfl
v3i+v6nzgOTH36LD6RkPVzPYT5p3CPotEzpYe1bXsBIjiMri0I/rMUFaUtqFheZ8
uQXKjbineVSRhgxml6By8Sg+g6N3656/FGTNIaHKU7h9irD8AuwVvGmX+QCcni5f
lG0Rb/qj+M71sudPNxG7J5HdiGcuyNw25+zkG+PMjdASh30HcBqdxDWt2k6VhKD+
0aOqTdtH1A68esRc2aqDt7SHAUp0skL52fi46EN2ZzKDH+Z+Um5YiFu8Tj6EybS3
l2pfFR/HPL7/rBzCs3Olqeql2K+dP9rIbVjKnv7XKj7bYi+jkt/RXO9Xqu1grZKG
gtLkv5/qGQM57L5z+1i46Ujo3t88qxa+Hp0kep8cXgHFZRCPDbs4wAlTEb3MNFdY
Sy++nTmAFKFLRSH0kImFySFHM2XBmRLlwez8QKXl/bn07ODJsKF8dqerhsag3Fv8
Oc/jXFKQk8M0u5sat5+3N1SC3nW5Qf85lGJK3lWprQJY0bIEC1oEn0wpTTbHFCXR
EETSQiVy87IDZMUPj98J1QBugrnVvtw+967Br8uoZYhemwIww/N+b3qKuALzyXYO
HXDvmYyUeDIMNreL8nFRvroe8hZbAdRxDvn3rU9yxbnoCw815O0O/tXbsguF4+UM
iOK3OGcNJhvHfXhJzCfsz3U51I08PuP0sRXwupp8LzsgaIkYocBsPnrSOpNmiK4N
S1sEIT0awuRQ9ZXytsTqjkJ48ehN8u0ohKhsvqYCBJbgL76nZ1h0INlSikTIAvyD
BQK1fhWYqxJWks92PM+kHkJZ20lJVNPC1wt48L2MmgRAiIxSVJMi/VqwoRJ/8x6a
SHmhFWXNypew3c40VkuVEL1fpOkcS5+05xuLTqeqJDKNNR1mf/LKCIiTjKsWfpJg
lRkn6ODtEptNlTKIVkkJjsIBTuidnLZLHykZC5vf+TsdqgamzVCW+EqFXejZEB4N
/DY4BJE/mc2VXvciF/wOOtvCpaMFnwJMGhMNePZDfnQJLKPdj1lREXyYfWm9JChF
YdzEF0O0L+/FhoMNUXj2FxA9v5NP0VGXcIAkjZZ9WPv9IVQBnAQLXAWmplwfyk4D
/vCk1elMQi5ZfFb16v5zpgULGRQQR/tIhphaxNPAme/h0NfdshRAh3XyRoXONmis
hturoj8uP6gnYi2e1R08D9JvmQ7jP3cg0iFUaR1Ejcgz2ujWmXY5uWbJFCIZXoM8
/rAd/KXfohDjzl2/pSLiRdr1qrgwUVTaTohB3KQiTqGUJloGIEK3kzPlLar7Rmx+
/xj9rZy2QBewZtjgk+xCzCcmf1JhxW/WyTsbTx44k63oBSSOWBvyE8iaK22HsYh4
TVEo2/DRq6sZhJkGLG8kffTHH79oz/BJg0NPTO6NnH4CsrI7Pi86GFVm/6muabAv
K4wdtsaNLkKwkfTF2Uuf0XZopi1KQttXfWEKtI7F3YUNh5ndNC+mlo0NudIsZF8/
QpPUmP95UO+Xr7sLl4ULs7jEENCRvnw6oTaKg9LiPjcuV2oCYVFLSjVvvS7epbds
2lyBmPrv+CWfhSQWq6fPrf7dAlMPSimDbln7SaOT5LgGaaEEm8jVzf8K8Amzq7jN
9leuD/DOPG8WdKrMG1kHXR5WRa5GM3V5j6qKNN9FBLJE4jNUtY/Vh/sPkDIjvlaT
hwtQyDVh3QTpLIpdinaWwBgP/a2/i2R29pkA0ynshVDPk+Meq48IZ28MUp96ONx/
/OWgeZIkWKatmPQdGLKAc8aY4aeUrsZ+cv7VbrjzhDh6GVR1YmBNbEO5hYmoELSt
DAwo5F+sKbmwRlOv0+nCQk/vJEU8BBd4VfKgXlLlN4GnMwxDvhrWUX9wf9End+RR
Ri+3vAD2s9lfC3iOVLeS/XodERwzUCorpTD64GC2oC9WRGLlHsfb4LgKkhUznURW
R3geLBxAV0ozLGTyz9/mvn98oqPIoZq9VbXxgm4miCwlkpBfoJJlHZ33Pg00c5Zj
b82bo1xiVo5dNWEri5TzdG1rENjypJc57mHT2le9uYCTntIhWqsvkFfQeib/ljpi
odW8P9MEMc19NX15Jia1yYeTNt/9K39vWJO9lBam4jTrT0xuDnx5rq5BuWHyWzts
oF4qSm0B5ZGCBnYM2dwmhI5prvyChf6cDtNO3I9xBmK12iLv2zZNgLQM+fmvuTBO
YuacS80H2KFCWXSmseoaxHrCrZi2J7lhRFKxipiviV7OKEKlnu1efXFVp1ScWFhJ
oEDcdleae/qPTVyYrZGbHLT5XrEbQJ/tQGTnX96FiUxzjZtMH30jQrEm3dhxFNj1
S8YG+WoEJ6J5LYRIGpWFlogSG32g/bACsV8evbTsO2rCgHA2TINsRBHEp13yTkPz
8kJuiphZjhcuKh7Vd4jiZWRQXKQHOwvPFcW6LvfgyrYWZqtkBIpFnoOWTto6NANo
DM0ZIAZimF6xGsyVTDClbwqtQD9Jd68Wsnz6NqS1ZkA1gtOOPuHKgWa0SAV8o5gU
PCRlLYswuqxE6IUeF2cvDSwN0CNYPbZQT6oSq/edPWC22M9lPz9qUR0D18VoOw0I
lx5/PrtjlUzgL8OpWxO6iukKMibHKn9q4699wMKi1AW3miKNh4B3mMywOKG4kuKg
ZA6AKmpAZfjsn7mASa3nNEnw6ycbC6myjWRs8p9lqIGG1ASp7FV6PTZ3m6idIQNB
jt7byGR6aSVxg6bFGywys31IcDTRGwqR1b/bP5t41nVVzq/naga/M8R0olV9eZJf
Ttcprb3QlJwLbF9TNrR4fpvnpnKfCe6vPwmpCvqP1igQVE7WMIlo+dMyLDZSAxFz
8Ljz+qimqY0UFKBcKDuE5eNHHawiJW7eDK3qYgooDkXAv4OkxwcijeY+98syu8+d
qJP3QTYmPLqChDt+jbHJB+ZzFzOw6mug5k72ETKtidQkYPolm5i1TtOMJUSx1XXP
S8ZpgLeU4RTkC41RrdCR31QjIfW8BYbZumuo4gJuDxuJ6t94YDX1L59yXsq2oMd9
oLoQyZ0P6EwqejKn1SMQl0hQxHSMbJg3ufRyZ9BUkhWt46cgLbqH2nED24c90hZI
wiSP73/boT+ggxi6LMUl5nG++4U70XQ4T5gwM7iJNH9pgOL3lprh696wo7Wp84zz
35SWFpHmD1jgcTs+fjVRINZrKQmuPkW/RGyeQgXAIEj9hq2KaIDByjN/HNGL/+57
2a8pRLR3l/HK/8w+FE/6Ti4HPUQtjrKh/Hp8ZS97apH6mn/4lWziSW1aZzpBTRM4
soxymqZygge905inPcqlJp6Fh3C6OIxUg0dsnkjTkF5SR6xGlZMyZX0oROLDIoNV
JdVp1fG9d0cPLct4mwi2btHHtq8GssSvMFXj90aE5C1CBZgf31YTpDm5AEBYzXKJ
X4zfIaaM51vLduFehcQaCPVjjlVCkxdG+PfYzQJtSCuEyyxBEkkSBBAieGX4Qk4U
JeV5f2lNKMMeALANUE/Ld5uqSqaPfZOoU3h/r71Sy1jeYrne6Ks3S3k4WpBB9IFd
+2FjyTMeKmA6hWgBUtH3XUniVO5O0oVPFmDXeXP3DLtK/3bH/12iDev63vYYjags
9wFfHi2xCKTXBwBO+P1PCzliEUtSR3/5TFypPEmh6EX1ufc2QcpL7ygEKfOt7sWo
7yvY1CCOWpXWb+u1COsR1uwyYS+jNLjDwX0Ea2zHwGck19cvNdFpFnxx72pKXOyd
88UjT8ctxa6s4MaWubNo5FJZkjJgYD4tSHyhu+t41bnDxbw4dCVhvRSQ6kZJjPRE
1x0kwgP+sE7bCOHQYm51McbtSKTKlURssSWcFtv3Ys4NdQ9IcD8SK0ufVEaHzbxg
Dr4F/iBpNOjkYibFWgWNlywqfjlD6yB0zMD4Ta7bW505ifXj82nwRCKsWVLgTtrO
+DUzsUKZiROb53O2q4nVk5lYXIdJp9HtlN26mhjXwATJUU8slidDFM4UZCpkUOx3
Hi42Pb81ILnq4vmAvaj7SKhRKZU0IRkFQzQ12Bcxp3FVeGP26cVPMJLTNdRTT15Q
EWQoW3VPpJSelWVbq5ykIJNjLBSasy4qOAyGPKeUoQyWTUUcfNwRDljFb9L41H2C
LYnpj47DGqxBdDN+FFetWPcMxoGOXjjTsKFj+EDcK1CshZNBENAdsyS+WNFiHHSO
Vth6lnp6+Hp9c7xBR0pf7Edg5urx2rWPDJ+pHZ7TYn4vR27Lk6wvIyLrPqU8ITud
6zm45+RWjOQzsF6lQJimqV6k7Qp78mnSJ6vjF+dM2mFsAhoXMchNnpnRXR0peykK
ZZDctOJQaSrJCd8UV9mrUuP8hzfVIImOBE8Wteqs/WASAeUoXj2r9Ut9YWeu+yN3
EHHIhDpu5rhmYkrJGya93UrSWDY0dcw3HrwkbhfP43AWdrwhyKO1BxwvKC3/kqEn
3vOcEOOoa2psUE3/Jjcli731lYS4pu7JZtLl2xhjZpQAskq2xCjkJjM/s8CyQsoW
RWP7FP2QR9juVf4MnN6esQUlbe5YiizlAERtifC/OHfEdv+9X+b4TloltLKSyaUd
8s3vOYG8k6fdMwRgAPwDAez7ucGx8fw+q5s37vxUyq2V+TjMLZSjkYMGtrp22if0
IdfMzetreS0qaQXl2jiMtKUdbumyjUxBdxQS56YnpvWMR6nBjcskF6SviF1ONOBP
Pf+hwOw4nwGqN+ue1xriCZJUxDJN22LTzWeIlW2P45/Pe60rUxDvbK4dSc0WwYBw
kddI6kV51KFmmqb12Hv6bENfrBoSj851c75UJYNTUlawxoLOhyAQHQ4BRD3+qF+k
Qrytl1U2DkwXROkXpmLznzStYYQLYcQhEcomNCSBm1WJNtZ7kG4FhEtdHeevOOlG
7zcIDuUs7FBDsedx5HfPbip0hmwdNBL0UxHXlk08ZZfftfVvUVbV5lIZmChgtL44
SvtJgJA09f04gDF9IWhalae3c+KjpaUDpdsH8jDbTm1T7p4ZfeS2ZoyjNiYm6vOj
YK3waVdyQTR8nRfJQDnJp5WAk8ivBHwlxcSWIRy2po7SqvTFnMmmf1LeB37QdERP
1do+Xvmm9fLFKWAjvIJW2DM+F4J1mwWuBfDrTrskU1R38JLTUi/VlzDjfpoO/aV1
XaZSyugaJnbxGmh+PseJye9YD63cvTU+NB9YkF3UeZ7gfyMM4O2XKx/qL3wVL7P6
+O77I0e+vn40FHHklO8Rw1LtZp3UDvMnq6QpJE7FctYl87h+8J73X+jmgy7U+75L
SgO6oLfvz0pcUXM5RsKvYuoF691nbSnrKTza0JMI/YzjvPfA5Kc5CwoPUUVnQp/h
ZWrbfs8pmymUjh7doIScdAXDvbNNvN1r/zjrQUpeEuv6IqgCOUGeum/LNenZs1M9
nXclPAyuM+L8Ci3IAvOqZ3VQT0akuBt4RjLR+NhbgVix0Zsgw5mLB5QDI3CXp0oA
2VD0DtGkdadm2xDHQ/bSi3Wr20Api6qB8/pRgJw/yYB8o/DELM1ukmeUZKTmpV0p
ylMNTMT7ih5ggsImJ6MofV2YLa+6eTrC8N3noh6Syyt/kVYuoxgiHUYhM9/uOu0p
OC9du94ctMIKU9/kDIfmC68BNoIJNoGajKcuNTJtME1rZarsoXPzNTWb0N9AAdAG
rVoVPKOIg65K+Sj4+5NeYoF9vekh2e1EJJR8Q16oa+isUcwp3qMC4n8jfxVl7EyX
4TeHYjgfC1qKjt4NIAj+tCdD3DnKLTv6aPokmfluTOmBFYfbvoyWJ0qxbLns68GG
rqV3eJ9dzQnsPqq8tIGq2fYV8S8gB/F857KpGWg4im8fCS/pZG4dEYHBMapQG5cW
ODUH3MBLrPplEe7btYgP+jGw//2FRTmo7JoSzmperKWuQIzNuR3n6WDHxFxljb+T
LMHsyaxq6BnM0u1/zgj9q9ifkYtqvFyOpFRLTV2q8f2L9hdKi+cvgOEQZfoZzkIc
HIlFDr+UY8YR83b4O5DZxTcKhRgJff+4LiRjsRw9hjVb4/j6VI8VmsxysYOwxgO5
i/zI5VefIVZq54o70JwWBykC1b3nRk0FIAeteYNT90PwQ/D2DRS+liCawby3dFCs
Lm/+LT4mKy6sJOFyMaCMulbjqt0rq0AsyKv1jl3T7FDcmO8OacdQeq1rqlAfUMyh
Sh+1MRU/GDfoxTN8f3+9yS1zZ/qQu3reMJgTOGImifvfWq5kj0C8UxFTaQbrY+1+
hza7xUiHyj6yxb2Pcf8hp+fHxYvvNS3RSOGxzDaQVx99xHW9CzLh/Rf7nKiebTDA
+NeObM4msCfVB/Nkv1dkhd/7tBkAIGRJU1HhPyC87yIUE44rIDImvd9dWpmK+jgU
TW26ir3CYDenaTA7Dobdhqk2aO8/oUxRIERYSSz/ZVVsXXtuvZGlDuO3xtKdObNK
EpZGiQbJZRwqtkjIUutaVnT35cLWReH9A7FJGax2MsBIyUWg6hjyqlnx6rTIYBD3
CRiqa9eD8PYxKIg5FjNaWrWEyXtnQaUhbxHHMoh7J2GP5BsliSga3fEnFitDEqt9
epgRB9ZUttS/dDT4Y7rYkRsj0SG0Vp5YWPlrxhmwnq7Y6ZkkU9C6XKr3FjMxrn2m
FgDLAmZjzqhV8w+xR2A+FnIqpkmXNnjO1Stdc/Ht4dqkualFOAXlB8FZJ4oHlu00
jMxqpDHRHEteDPKx4Ux8ohKWvtNY6ucQ+Hm8g1TOGg7+f07xiz4X1VlJ1/2gmXS9
a+DJEwSscHyjnot+6tAU+HpNwaMUic9sA6iXqqgXC8yaQF7K4lGVGF2HLv2+XvBz
JbOu9VBAK6UohzGqOorBGLC/AsvLsp1q14drBVGS35Qxd4r5CKTM3TRLOvN2wTaD
QHlUX/DtM/np2jNDRja5yuPLw7AI8546AB10XZ5noSSvR0v4DGPYkr2/Qdgl62dy
4uKdI2s+NxQDZLtT/JPTlW65gntzxt5AM9TVxRWqKlaitki9RDRxuBNqBbTdLWP2
xxcaH+dm0gkS2fNF3mDnahGDoJPX3ejIopHhLWLczeI89ZA00LEvyjKV/P05vl5g
uZ4hqtOnVTJhVBO1g9GOYbe5+3Mnm0FRkmnoZwekz+RCAhkm8ckuVH1zpXXDT/GA
Uh6we3ZsKQgCCfrjmCj/Ba0U/n9tJjwiSg9mqs6CiY9nYMR+LObhq0070Ir/AoTZ
GVRhFdFViqJJHCmh9EoOH7cISKsOJCQtZY1Ot77h3JNmY+L2AlxCSdn5c99K/W0m
eX4xBx1VFfaTH3AiV+jnzuOxcSyCeC+KK1iDID8bIIvinOmzpaUE+Iz/nsr3KJ3+
DFRQnINAMJJFyFKe+DAb4UiGTY7tZvYKB0cmXWCVJUK7aC6uC1UlZIrcwazLfXjM
/lMIYMH77B4vl067NGcpg1w7lJM2kj5BFYGPl9r0Dh6NBAap+0qRSlG4QxpPBMqf
W0BYKclGQOuHNfpMeA6SokJJ2faBvWJBX747B/FGnKltKX98ieJ3D/dFO5m9EcOs
oiYTyVUwpoHIvmOdBDxuvmFcz8YwWkDjcwwQCDH1QUvgz7u1aJ41eN4BwYGDDpug
t4tDaBCi6YLcvuMg6r8LZtNY4KUgqwnZ6Jhn1CBRfEKBGUeF3x270wNzm9mT9t9v
KLfZE8v2OiZIwIvOkjhjPlFDAAXDgS4KhLj8XQ+fH7MWagXS1U/vV8N6B5NFmGDU
NuEEoF5402ZbVaVxLeY6t4gh32Q+P3PkxH1mRD2xob8jPniJ31uZY8IqKctIPNHM
ZWKJ/ZUR399cg03GVYLe+bIpJppxOEJPRMueuanuALFDdFslkaxyGTAdQ40C78lr
QP8ig2pTLVJaE5DWdQpMiEOwPrG1wYDZZB7o1Aiu2rF5Wyl6+gpUVuoiBfuVBlcx
EUr5CBHTCC+4XzeZw2CPHUAMYuidDE8sU8r3Ni9b4I26bWHV4dn4MXsgug72RU3g
GATMZJfqNIN/7SAUCHhLJ14n6n6r1q9vcDpmZSUD+oDBX5LQVIB65tWXYTrhajQI
P5QSZP5ARXhX2PjeMHg+q0s8vWlxpkG/1AMQAX+Q4a+3VG4nrKbI7GQ2FhBu5xI+
tPlk4JLtMXTgKmbvVZH3Rmdck/urJTqPZaO/5lTVuzGWjvHh+qvLgkAhHldLbO8m
Ukr8jvEHHhKy9FUAYCbLHWRfYWePUnn3xHDEYMmmizVELMWYEhHp9ph6e737ulXI
GPUmFlkEfMgnkaBx4AKJh4tKB+yoCREJWnjOUGLvVQov0SdQY32RDF8XUtYoCTwu
6mY0heidrrl2OFIoVXzmYA6Jh2FsFjTO055QjSxTUfbMR4ktz8Yukdm9HGQHqUnH
ZSR6xkzHVc5cKY99xsdHjz1ztHlZ0yNt7s2pA/aFlUCj89uMil0Z2sF6QEz501Nf
3ICBjpUC2NUhA9t7xS5mFIG52gKF9bnKDozruTHoHSSmp65LhRYUJDW47Wqy5MoK
2uct9eN3L5TokvYnz2WscGwcZf9J5hZNrTXYPL1nOv0pLNElT9/ISE57OvXYXrb7
Fv795gPOO2TAwp9mm+YCo6qT52NN25rsrMkwarE0EHY1341Z/2it0VB7QdWeJmlh
p5KDrTSF5Kt80wKZihBCCDqRmvXO5DZMHEfmgB2e9EmPEpx553OzOro7qOVjjZqC
68lpHLvljf9rslym28AeY5VUFsdFCigEI/FC7EeUWyz+5W2xWU6/Eq9r1NKWBDpU
4H2KjoVYrFytBaoxRonqzm0uQ+GRXS9x5Eu9R86A4jYwGrrc3EXnQBKVESolemXC
Sodh9jTxW77FNgWFKwaPjau/rv7RYGBZdbZn+M8HtK+tS64SjKArXSYXMELoSMJS
uG8j4kdDjLe5XEO0O3NXtCDqryVC7TV6y0k88PmMoOMPHOPhtjHpqRf05INrLDuv
Wj/O+Tdc/gA5636hTuioqsMjLzJI+bM4UStwjdPAWAGWdf1tBFO/RJ+PlvNfW5kO
tC0NXlOHTAPwbMin68ugcTy6Tb+gsMHoahhaTcTWqR2vgg+j/RslzRHNw2SpF/pZ
CiMZ0GoIGB+gYCdduOewYXq9lShJ4bIny8VoAGPzLrJp+C7K9o36vJ1+u25l9AR1
+pQMZF522yjHPiCWr0tQv5U9aBSIUulQePXH+bgGIWLj5UCey8CWUkl+fvvTVyjh
REd1v/ZyD0vTRaOzIBhvbMdPz9wTYafuvORbsJXFAJbKIZff0QVCWSBcjhb6H9pt
lXucioAx49AgwHFD2v0JeRJkW3JMx7QKdbH1rN/mBiIx46oHXZM63vDkYjcQzO4j
Xvp8P5YfX3dj/AGL5/MIz4YaSSp04az7D6BizoyEqqxuyjDbKwgdfXmgHiumUTLN
Ag9FCsYIZZc5RS9JzAYxkBRvn8wJuxP9FgMwf1R7kb9MuUPoyffzohDmCUllGh4Y
IqGr+i2iIAsdak9faA2UseK5z3GvSfNbaStE5R6yNlf0/V3dTmUBzZ+gLOhNuEZV
G+oM7F/fpjfO1cVtnHYEVmEZB/RRLWia76o84wRRZuIp5d1rv/V7u/A4HnIHN3BE
LFwaShazCAjme+vNVRx2hfovuzJhb69ln7HlsOFz+vTsMQ1xbbmIhArkfE87yjyX
mYF+OgyZSPQtOsf5dBHhSWXsS53i8M89Ks0uOM59k7bhaSXyGxVxb8WPZoI7Ol2G
O7TwSF1fFLJq/7avTX5OLlT5E3nrhPNoOxhPm1Ojq+ZSgpMibqJIBxDPDJCCATJ0
0hM4XLnqGAeuPxqe0KRjelXrOu82c99vB4FqzJrENlu0fujMs4CSM2gxkDiYT9Uc
t5/3tLYdm0NXIaXuD6hrRfWFL++hTCjqoO8Nuu+HkR2VdNSVvVHcbdt1qOS7/LmF
Xs9v1tvx/1oR7PPrqXlpxZ2+41LXJRMDshBG7LIW09w1bl487YUlRrY5ZSBtUOyK
H/sz1LAKUaLYugYAd/qcHO4+Sm6ZUIG3PRmTIpHGIwCQchP9sZ9WxgeX3RdslL1F
AmOwfzN7opDB9HsKrMUCrk3P6xDjuZ5OdVO0B0y//abBweoLM+ENZeFzWor8TS6i
Bn2HFEXMBsO1BfaVk9/WKg3/1q16rCUkOk3Wn0ERQezqURexm/nEPQc3/rNlPwcJ
a/eGF+R7xoCaHIS/dU+hbt285rjPOIy8MoY7DafxjYJElc7yDz2ybO7tO7x7VkAL
2R8Q8PSfsp7XKz+rDu1HB81lDPz53kCDbQde6dtiGzfsOEX6s8GEYpxZS+xweXED
dxaVVepxrKfOn2F3OwaO/dSOao96DyPpVW1lLJ3MVHbnyeHpj4cJ4/1vfruPanDR
D/PwDgmwssxJN0rsOBaTQ4fkte7wSvw6H3lJBh745y7BLm6DbFJsCXVh8QTJwess
ceMCmlwt2RttX4d9DNgS7CdFY5sINzSayd1NL9siaJ0jtFT2LMGHeAfgwoYBFf5H
fkJ3VwDArdUAdngeWt/Zaw16z3ho37FOyYTi108kP4OPPhWr+ZwwmdmNPYNxxBOh
2yM0TP4ZTOX4caf3fQPCIGLh8UmuQ8JyeqKJkRLtalXM6ZIv3xV7lwf8Oh4rKWQj
ibWKdpBUYeaDwMv9KzEhz+C8VZkBSpqNBg4YzfZwjHc0EEaeBYAqBmI2vvmdxOot
TjE74kiMbyl0LDgNqfk66E/F1aeXKnsJ4NW8uMWulhwLoQqmS3bxSskx3/Odtmp+
iO8FoXGND9iWwztkFmXUar55utUdsBKgtB0/30XnXsDbaYqoz/mXSwUM8CdwTclk
mVflDiXBd0ymBPb6n0Xa+bvdtjCYSHYyYsVO/mK+7PSjxCfBDFukXtrS5JPcUYsm
e9C4ChRbn1G+xVdXvaN8oTfwHHSiusKlHFTnbX+az28L/C8f0JOj0t97o+ZJoxXD
T/Jci4u2evpaomBSE48/tSIbNY5jrlpxCjlFacdzz0gZEOlrEDfWEeK2J1gfM2tF
zhgBHuUyKDUdc2JMuze75YXzi71mpp3dV9V8R+kf229SxSNIuEA8eTt6ctLfz7PQ
d8l3C6gXr2CUVZU6u9f34F8i6xs+wNOKBEk4bgU5K2WMsTgSgehpKIjqvWv733nH
S8o1MSUCSl/rIPsoIMeAXSkGa2hJj+klb85kf/p76Xv+Rhbj0QFvYonTsMHRkChk
DVTH4f/I7CLUg+I8fORkrLg0s7kcBCCFWEVvykz5Jk3FzoRbVXFzUNtsOBBUu2Kx
MXSgFCZoev8BLismrLuzx7Q2VQ6J5Zk5KroglnJ9AwgDwcA1aV5asIKuMeJEZADr
EDlDhpPFnxZIviqladDvwovK1Az/mn7nK4CHpnYeMn88dlUFw6pkzOtr8DsAPGD3
LcVsK40KPkbUMIoRdMrHsL9ntBbwiNyhpc/Kqc8EN3pPOrag82fZNtvmPCCJEyFm
0PfD6GKcxP5ZzGI7HDdFCIJnshTFZAV6bpKmFpGUP2BpBTE8yIL65p+tid8etMDj
o5UJJ1WJ/8H/TJEb04txnkoL9NOyL8m05vvJx3ifaVKHWiOm8zj7tCAFkiaew8a/
kC1gGlz3ksGaUY45tzfQ1WV4eOCtjYiZUitktrrRh0yJaV+f8uY5e/0WuxVFxs4X
XSHKovdB64WtSyaj+FaBesVu3ylvXYuz/U1Qcrl/ZmxuVfbHEkBAbfxjxdRIv3E5
srZ+sSNLokxaMaFh5na/MEmVAXrxu0zuN/GdpO6m/5bbHCjEM7VrdQ1FA+yHkgBS
GaBEV5mFx9zAS75Sp6m2aLS6N5Xm/U+vEBDBb8ggQ2C95pgZ9dAFWOprozc5CH4X
Do3g8dtfsS6OBdS82Z8O3b4g8Scns3SSzQ2ieq5JHc49xL5jPLoz13MPT9xsVqy5
AeaI7QG+wPzM4EPQJuB5f5x8rr7EuIw0lbH42kIiP4S8VIObrYtuw1nVB1kbjr1v
3DyvybrgMWmNGk4c6IJ+ucBva7hUyI6VoPM/uaEzJZ0kF3yyr2kDthy7bnnKIBua
TiAd7+qJDnsABGDCcJBmQGjEzJ22i+/02VQolHIgqf8JAUSjzt5CIswJuhJ5A0kJ
2MzMyAnfInIEfKrLCAVSrbDSU3zISgckj9FtN2Taz29Am9WXLZwp/QfaKmlQHYXP
v4RHi5tKR/nC4Lz4tZaKGoulutzM0cKZq0WC27QtNfK/qqoGxdWBR8mtATFClXx8
GGqQshnqpA6iRkfRKA1yqBjKh6ZcezhwAf1OU3370HXjUNY+EQlVxZk6v7fDg525
FL3vCOVotMKxzwIk1G271fqJPYgGc/SkCsT0vb0kPuF49zUq2hG8FT4W9svXDfWi
dCirpnmKk0eM54NKk+loQQU4pwT6sBxF6JdsbeXk8snbBHUvpOq63EX9VvoBuh4p
C4TwKjwQKh1WkwQDbYLFatsNwCy/b8UerhtEO02Hvk3rPw51JM6oFoDu7G+uT0ss
YF8mSupROAQZATvbs1u+OUXw9BCaF2H7yLuGFViX9dUiKaSqQTaJnURyqJbSIb+e
6lATebndpUwpmug5gdIw1ZYo2gwIZDJWvCWKE9QNlA72aTuIdkIesE8WD5gpGNX1
TqUNKM27oLFNbShU738NnUtHBM4gUbOiGUQ438/4IgF4hrGczVlUFBwaioxzZqRB
czIlXsdqJK7qzQitSNQJslxBmRE26I+5KI6xmOTGtD3Cbc5tRo4SiQ4uirkFKCSG
z28M5vAUtCZW/azW0Q8pCvZtugDQpTeWkRb2s3RdRYS8rQ1N6ox++bSiG0uJVZ55
VONPSeLh43K/QoZtgH8n6OiXbwzYDaiUZDSXrocbDJThgKnWdhOjQHxYiqdsZCP5
8KnV7Y42jtCiPKC/y44Pbj7C/fHzczEtkIXnRxJJqtUWNlBl6x50f0cGMrzdWsRo
mjFQFT6YSFVUvv5c1Kbhx8cpzY5fgi/qd2w5nyALrlxh37BmcfVnC+M47p2I5H/9
io3wpvyCy4SkTsnf5GmNopB8wywm6n1vnAySGIzLzj6e1rKaOXvXaYCRaFLD0XfE
pVzhsd2GE4Q7dZtao57GN09apQDIef9reDan/lrrZsw9/62AioltRzzoJ2zDcary
/pbhIwMqld9lsHN4GLik50QIafE0/pl6eknz1hPuA93ZNPzwqP4T0CTkROCkIXO8
A7a0Oq/ef6w3MIJrsvDZ54ePMDgwqoG6HFgyQTE/eAnR7psELlI8Sa+gFJJwUQwq
LtwDkjP2wCfMxUHQ4dlXKbxJoNp0ofrG2jkHEzDPuYlh5OEIQLwThAzbPHKCEvpd
uZZNWR48dHL7c38ikBO7gOcloSRrICTARQhQbmH7nEU2DhWItfuMBWQloYW7h5uX
XzZYmLw4YBTZwMo5K2rYURgKZ1Iv4CxFItXMoAK0Tm2CVHhV2KhBYYH7DvHma5s9
94OF6XQ/ZVw8AEzO3FxBxwS03f5dRgI8zWf7xzHXuKldXsl2P0SfeYZ619AYVilt
eoE4g4mFtj2V/bqqMcg7kXU3xhaTvwA0t4KpbcbV6pIj5XRv/TJMtDQUhX8Rj/5T
0bBoHyw+eT1Ldy9sTrhGs33KR79yenqEUTnQwdDNrT67uw5grI//JnehlgW4VPUL
pH1D6zstle+Dc3c6R4/CtFN5JJ4IKqF/LAti9Y5KpJHwny+hZHBS2Cwr7M8pRD9D
kqa9Q8wQImzHf2iMlnArIJCKb7nzFxoipwQOiOGItXCyI/bCmadeZOEu0IPqpCxe
jpek09r6qkO1MB8c0zMJ7wSNS37JtkMlDh+zqdOtTLAZnT7oN9502uq3JWJI5xMA
8hYF4EZoNpyl114JUDZED6l8zJqMcag3twxJLD/UsJtH467XXK78xP3o5heux4z/
Q9Y6WVYyoXjCOeQ1vGUuxqrhycI3JtIZs25LJooNCXnF7oLpeazZPWeLtnj3tv1+
OS2xbA/XZcpHmpPurQGfRDA75ao86+kzp4sBP0S6kXFhCEsIF8vqFLOMiREUScav
lyEZSBgBOzICR9Jjzz1zkuJxa2c6J5x+ERwLCK/j16XyUmFHew5jGfwYvHpxS8YG
RCWxI6SofWmxyFezqt4WVQNOr/4MezTyZ5OLI+Dqptyztjx3rbs0ReIuNzQmE7Ef
MovMC9kgs18gXrARdSuMxRu9H/GFBNX0+se9kwpfcXdXtpBbcyUSxTswdI4VabeP
96Aj+6YLsYYUp2Ug05RFoLIdYhEeQ7XRBc8gENn3NIo7ju/CqdB/iR2Hgb1nXKBw
l66lcTgH5lbwZKOwasgH9j/ra4DM4TLI/aebljHFoQ8kPJ01GPYFH8C/5+Yf0kcN
2e/zXtq402IUcx6mm69F33toSj/NkHznFMQCXEdWpS8qAgYiQJO02ysXnMwtmckf
Akuw1EaVz6WAArpPdMRCOxt/2qq884j3SfGgjixqm1aYZLUFP25MYtNXKuL0Fjhd
D1KrRZUwCV8zVuZbKS3/1Smcmv321gZAew4JVuph1fzbihK2yvPy79g0U+c1CT2V
lNRfECWSU9iXIYNQ91Trz2w5TTMVSflMkETsWq8RPZFO6yy5yKXxIYF1ukb3lHcI
bTZAt8CKxYrqsN0l84SXi0Nb+nH4M/w9vdfSg1pN8Ta9+mEsDvPjQClu67dhXgLw
PGtOdDL1t2ZFqefMjzzJhWXwwRCZQWEn2E8kA4vvWTJ64DDkZrkYY0dSq/Gkzfn1
lAsrWeODpo5T0x2TastHQS4QbkXJ/GqVcmu67iYwMxXXNXx6DgxRraTPPj7jRGV+
rAWZIktVUxTRLxJYG8S6FE8qqabpVIQZ9QhCkjLKoa8Pr/YebxW16tbTCKmTtsTP
EIbr2tukEUnrSl2Qhoi6zj+bFcmwDivxJHv0+f27OEoPuW4jLYNncqClJBiKdFSq
wNbgG7v5SuknEwhLwJ+d6gTh+/GF4mDo8AJibgwgVKqazhLb61max4LXRuwm3Xqg
vWMeJi/N3L0Bkk4Kh2QQOIhPpuy4kjFjXxGrG6PLviaFVZHItHzlkLu8+ym60d9b
YxbTf5xkpZleLdlxaa/pv8/hOyehUYSPRQ/6B/LmjvAFXS9+KXf96abIivqLYFgX
kDMCnWG1yiziOstFTTP/3x7PrADatr7ff1Yyxu1PMJ9n8FuOhRu2tdvlPzD9oqeM
YUHyj85WpBbcEkoBu8a3jXGV0XurALLmwfjGh+Ha6aq37zJNa6ANhXOc6oW0Vdj5
mqm+uNJ4iNo9oArjorSJ+Z7ZI+rLpdmEvp0YF/vljOpGOSmCQRAGelJUPgTSRxHd
WP5R0EBbipxfgyteKyDoJ8DqQ/FPFukNmfZ+oCzMck1kmbFTiqmhQgLwvHdOwkuX
m6i+bkxFHTntFiGRLllspirVKg2Psc4TKhqb/5jT/dWB+lGaCyEjyicMwV+r2xaA
uIpluij5QHkH+G/u8Ub1na+U07IUjUb2Jy7alZ1BxerYxZEqgaLZFY1H7Rsb0pgr
je/zVflVdpjsi0izK9RkLVVwBwUpP61vGhLQNRa0Lsev8qTj/iH+yuiaHQ3D5Teb
jvPVNlsXl99bX3aUq1NMgiKeIwNbr/HC0ePTWeOulqQAWcRVC1fFyNqsstpThwPc
voX36p9z3sBuv1JOwrndXQCn4Ot+4IH1ACiIqPy0zYV65O4s6CpeG2IK6yQmLrWT
MiZsd+mtwrPZxMJ4en0D++/U6PhNz2Uxe1ww3Kx54wJ+rRDGtsobgNtcOJTbZ6T5
LKGjvjmKDFwZ0l3Q2Z44Oc4bL9O0WU74AlXraI3rXGVXVbXuF3rPCnA/AAxutAB3
wxmd2HkYBHHIDflFUbd8lSwQbsftgv3Bp/8cpVwb80sSlBxk59Cji2/Jl3nfBVq0
wGmV3YEn7DKIYDKMLzTh/2IFYxVuwFOz47LPqg9YosRMRqA9pYpyJhnVLLb5Dmxj
uuyKN7A3S9Aav1sD1PD4lJHpW6AH3SB4mg7YYGLTzxcPq7mHC0vhuZstlawXp7ys
AIX09CZAtnHGLj59aEW1amPXLV0ZwJg8asNVbTu6/5U/s0aHBUnFBurJiY/EjVO4
+lvJcGSMQNUBnwQHsLayxUXS7v+btw7miFLN+VI8nzI2QsQQ/YVWTRp8ZxBt8TxM
Y9iR+8X1dg/c1/wWAu7/xux/Um9Z2U7YKlSY5AS//IAFlrhj7JL8BcQV59pB/5cF
9e5IoJgxLkMMiO4uWA8Jk8WVTPIgLvwNCsZqfEL6kqblVoy4q6VPiLT3O6D3MMZH
aJtGXdVNjrGYbybfDxOdfn72pVE04ppLkf6rauhB7o8q1EUHZm5wC/geRA/wMV1X
v5+02rM2IqyQHQK/MI/BpACcEB7Jt+Rv03BRl6RDwCQ9iKN7rjh8eKUdDmdE1lNs
7DoKLWmfNJdBd0DyGUlhs4FZSB/3oLuUDESUUVNTCOuuhWc+XUKgawCCCz2PuFAI
nB236Br43oJaY/BXf6FUa2bmTRDCsKae6DNm2kVcZLuwSpo6sn/osHjT2WYgA7M9
gYmpFkwq49khba8KHodDEUaU9TlU5ooOYdZeiQuU/L0c7SsgkG9InCIJkTDUHN58
OJCtTrakawXyTmEzL00saULOHxVpdxYGj0iAiztk8Fp+DJ/Aotdfz+8K760M3xRE
/33mrSU2z+JJycrBfwIZR8SvSx457QO+eYR47JpMxnNrbFmQ7QfmxEEzp5rUqW9n
kREsvRMFoYw9S2l9+nPV+j88mXkOItpMXqlxvt1aC6IzTCByjpOqOlC5gmWqQyy9
bTVWtbcxYlYqRdGtOC+Ja1p01pfkuSuj9pZJHBURS9/yi1mbbtyweRv3U9aV9V+L
vju33xHs9J2Nzd0WkCBIMXRz2qwmrX19OxU8agmhdejBAjBbEUZyJAndtMgtY5XG
Vi3SESREyr29CJ2cXZAy5IZtVZfZBOyROh2Lx0Gavpc8in83bUuTaDb2m8E0Ht4k
FOuHOXNLFv9jGAib4/EQ/yYfE+I2Xhrke2dBJS9qw+JG7dyojHJNaDwXZl3RoTC/
0/NBE+NVGkRl2A6hdGmb5ScUV07Y1dfymJYRU30jIxLngIEAjAR0lp/ktNI5mOTt
WZxxz88TBGBp8GPQxym9zyApue0SoTlsh6LQowk6ydMmicRtr2BfDY6ujT8w6QTz
WeVGKjMoWxMsIPxnMRyI56A6zjvbme8AbunsWnvDLrPrIdOEJPHkj3/VT0Lw5dmp
9VM3RzKNgDGyis+LqpZajeM/zzDw/OQ/ISVjr+8qDsWuQeX3/ZtM+HfbOCgRId4h
Hf759bxziGNV4QEQccq7Gh/2A6e1nuQjYX6AybqJBht/bPTWLaLgZuFbZe7mN0b+
ai+fiI3sfurq3rvEMDFTYw83ehfindemDvhyi8OMby0OZnw0oeSyE7/RxaYoE6VL
2mFcopM2ckrxBqZSXjEk9pHuYJPnEehegM/Kai1UHBmw+Z5zydUvANz5JkD+fHYw
Jl6Pq6zk3uCPeqYQJ+gamaFK2jEhWqdkYXuf8teZ1+HyjBdoz4BGWxyibrsSd/Ch
ZpmXw1hnaTKu4m8HiNSdMmJc4Pgkoesw7C7dE+83KGZjq7jPTiuCI9d7+vbWv4cN
0NvTf8aVpZoKwdwqaq94edL2IyONpL2no4j0tUsX2HYvDSD/YthS4ifktRVzqd6w
t8Fa+XcLH2p/3B3XOSx6iIXxrcr2eOvShbH0YEbhISSu6BySsJtVnaZFCSUopTXr
UmMChp71r23c11dAi8hqYxtwz2/pJH4Q2rTJqYvQ8fGrtVGv/qdxMEUGYJaD02B3
9EWlXx9gfdPrKLqlAACAmxg8WIriXmPzaGGyZ8ejc22MumdNKkAg80ovIpOnE7vy
n+gd9KQGXYsno5rq/sk+8Hos35NRV45jQ+pmCIx9JO0vdKynRwh01T2+h8ye4Lbw
uwJkx3kVECpafMAStJcSXf/AoPIT11pG6bCWwrGkhyJMmK8w+/+DfKpdhbwHympD
B27bev3U5VeklSH3+r8Swfp8r8ddUn1oppwztrrARhQHxt8zYA/L4Xdp1gU9efH0
fhPNFDBHKbbFDzZCxrrAo4chvelFH+wiFshRL7AQFMdrUdRbyF7nwrH9Ml6qN2ot
YswcU1ecDz/q85KSjNAon3y8X60rEKNDjGJ7fUK7xqTOlZLcgjwMsuWXK4+gAsJ5
M+NFPIKQpQD9PS+XuGPoxHDz7pJ0XyZTaAWt4leauI0CNHf306sCvBaL7Y6vSEKe
weAkHFPS1xhgnBLAE9/F57j75n0OfbCKBVYOCdEKHZNY43WBOSigNvCJL4GoNDkw
E62bSvsZEqwZFeWn7RjRjG15CoKLSpFlNpXQU/ey278gBkM6ItCRqHUkg5e+AY8+
ztYWHuVMtQ3PuRKbNRUHD663KxwZcfE0VtM6vwyJjQetkCT6E38b1xA0DAbS1k1X
ISIJ8mRjYD0YyKWkXzNSyY+vu/l4ekIqA5ntH4IlJmxKVRGdgcbAEv0rop0j8Ctn
VbbAkI+k9LcOovRKO9RUZGsf9BdD6hU/kR4XP2072pn2ycf0zurgVqF+dVMwOwd6
YgZmerS3qMG5Bx6gJWaoKe68FK38CCtsMyfYsuUL/Td4PZDIR64CakhRVNh8lVJn
Y47zQhSk/+9oLcPMi/pGp5dBGztnIWDmZFicIjrt17yvWcIeTh5uk5L1k/cH89PV
88quNz/EXIcg88W2K31icboZ1z7HObi0Ap4kLkeulQDH+o6fbW8bBXIwHdaLHEF9
6SGtIFM9jY5S10+oHD+sK+IWnEEYWTl2i1rqsi3T4DcYdJW1cftzNaxxB2SgTUua
w/+pXwGpBdAHDnCHG35oerss0evjJ12eVDFxrOYSYNeykLce90A83THDWbeY+7Sw
kNJ/42QLN8gVVQ4WKzgyAhtuQYj6qmSEVf92IM3b2zvIKccRcXy+v0BPF7K2mt+O
t04xvFplTrRYpeyfSMFxn5XTpiYBqtE6pvujMXRAH2UBG9qFt3kDN1azdwxgRVPS
6AiUQjFViPN8kWDK+s0hptVm1A2jiVLqR1x6kM2bUrLSzzaK9fhA0OrM75oJ8LTR
InyqrGiBGlIDAnSxGWXSaePMjWiHKqCTkZV/3HGq4Ov0KkbHr2jcwQNwuChkkjv9
xFV+1BFx1PPTV46AuKFTV+MrJrz8kjihR611hEOvd/lM8WlVrRPk+tLw9Ma1xwWq
ynlqMzv7S5HE/0e5NFGfGv1tEYxey6GxwLFFRWiy2+mzgknvY5Oz2rndb+BXKE1A
aqVSW/o61+7b9ywI/fvBsRZCUKs++l/LvYq4w3eq1RwkvQXb6NXCv+XTBB6gbsfK
7Sk0rs9YXK7GNdR8tYxlhkV6DA1qd+FYssFoWIzlM+35sQFHf/VEvi+1YkgOo99b
oaBi/tDiUMexpKF5D2LIDesECfY1ZlgVu1TPHExh9cG2nSrYzEnRRjYKtODBsoaB
APz605hxTkAEvbUOrRKhu9pOyfDQVNjqBafuYmQUztzqLKPyOaRKmiLfcz/VLLCz
XkLq2mjZ1O8rGrj7GSh7t8eNVpkrt7CxUCwjNrLLOi8aM7yr+y1V652nbIQrd4fE
2ZJz5xm9AMdQCEjChUk+c85ybRDkKzWUeLsVKuyPh+q8FJuq3t4DVNaGPlTFRxvE
ehdVXWmys1KDqfxnjClApWdpwx3j4tdpZefU5RzVdxhS1kcE2Z+fXX1e6E50v8I2

//pragma protect end_data_block
//pragma protect digest_block
/kwGVy5i6NSFD8c3OtYm+SwUzg0=
//pragma protect end_digest_block
//pragma protect end_protected
