//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
rZoQsBU2TlF+3yF3CbKWgfrRaylj/p6aC8VxZHPtQla1CmyVekUD34L5AdU6l2bv
YAcLYe9RtCCaHTlRXyqZrlKCsHZMKFaAc9uiEGSnwsL+Z2HhUbZnsYIrXLneRmyi
i2JA8/nSPnAvUh7gjUk1Us14SM6hbDs8pzgzn+5dmEKJ4KJdbgDZKg==
//pragma protect end_key_block
//pragma protect digest_block
7VgcruTQGW0691JIa4mptnTTt7M=
//pragma protect end_digest_block
//pragma protect data_block
fHqJQiMyb6NzzWlIVQOTKi7u9ztDmSK0MU3Gt0Rt6J9ahUKQmU6r/OtlCzbWaEpx
lGI5l5HJCqKbD4A63knnIiu3uM30rLbtahg8a13dF2V4scoARvkRcNm6LdjO4rBm
EPX/pRV1OT6v1ec07G8gAHsitnQvyVh4o6Z51qzRtqTktXcZ3cxJMnHCqakYpGNm
G9tV5y8i12XnJx4laP/fg2qWONPhq5/Zn7n4CC7Otrdlku8fVZPjdXm4KS7SP9Eh
Gh7DIVvrTPIMKoVRXiMj27CmiWNZT8SrNnxryyTGpEFxijCAsLRs24GhFHfFAJTD
3xKBw+7VXow7Obyfq+c5C5QxPi6fzJWsQuVUJVZrK8pgTZTei5yodq+9ijf5cfUe
I9CAWDqcg6NfF2ZRj6+PtFKSJo6ZR+rPU+E/UA7lfFmA6jvbHZ1Bkd6ut5Ut3V2Q
2+8NE3pYuG5ebubbimEutW02zx3tdCtYCW7cysfGv2Dq4iOsx6/2jzDHs80BSwxw
vPLrf/eKeeant0K19Ei2Sg+oeVGez3fbPHGUQCG67GW1FiIodRsg2U39t7M1h5yJ
W/VqXMpZx+j9H9A9fI1KGbC1KwW7X2ddgKS2BNjlRvdz5xjErWPyP5j6lF3y1FGK
mrdKlNDberD6wD6Dh96mfYXnflMyQ3tLqT6doBbZxa6J7ul4uIkRc7Yc8GGpOJyW
QD47XzzIl/gQZE+9Kr13cpGcNSp5JGllnTFlUSjo//CCllcn4Go+K7404SchQFlO
XlY4N3QpN1o7E1Z9s5tvv1U6q3npQjaDmYH8ikkAXDlB5P2g5r4xsA+Z6MyYz3GL
l8oP0b1DmNmBh11utTYag+k8IE4CpiuHIJZkeuWJ+Ush31lLhr0R3MXpslBW6j5Z
NQyNBWl5ALnN9oLzcKDsSS+6TzyeFfaeOo07ZLPizUbeBwTOwChJgsP1w5Ybi2I3
LjECUltUsBJ1XOkjyaer4WZyFZOkw0KdpgVFLb3JUllSY0/G73iHg0kDtlZYGA9y
VOAL+jbU9g+OIYzYRKkphQbAl82meP6WyW2gr/D/BEDUIccQKjmkBjYsoyec5tAD
pGSb5WfsHkexWgCOm6pd5KU/HjnkeQ3zTnoVceypvWfeTmhIci5jkb+lbzVmSbg2
BNnD0aQCvRCwRqfvWXG3zh1OSw1lKOXd5YU5/pKTbxk/MW3rD2pK6UX6TfFOCrEf
qErEi/FTxz1Ut4lhnRvVqO0hN50HCOZGKupR7H2K0SBaicOYw0504UZcBHpWMX1G
rM4c6KVCLuMHuuTFNbp2j/Y6OhrG1z41ug8k2WZHApEgCyYkzspzycRCEE+FklV3
vSsvPztjn6c0jqmDUhZDS6OUTfv3z8lT0uRmsqykTifFwO5M64oTJIVFWHwCvUvf
eGehAmmGKyr4+OM/ExwCqEeJmiRyEfb4hMErxmfudEmlGUAmu4dwH4lDEJYItZXJ
EE93gfNjFBKw1G99r3ir5ENtOOIaEY4eAf9vcHqYuXDU5Q84m0diYAFlQTVnj9h8
1F8qJPLDRcRFhzWlemu+W7lN5AjkWqltCLQK7d6SeLz9me9K5UdpKA1hn3Q8WNJL
PEYhU2RwLy3o/6DLaJRuJfVbe9RIGZzN4K4ti48RxitBAlGSL83E83p5kBAyHJAK
cHV4OKXz3zVhfGYUNxQ34SQo2WZOu+wFK13TDqEKXI3k0vMD+xZ5KALsTI6hlyxV
coGJp84TnvSbDwDkmuJgily+3vwY2LzVgY8MDulEFEaQYFIf/7RKvEO4dJtl2aoU
eeuhzw0GCpQoFENzS5Ew2CCXIa1KKOyt90Hv99k4k5ls+Cqgc/6qJ2Q2SFPbwGyS
uN4iEIzEgj/f2wihBBvW2T024jk1lDhaa2vov47uM8l23SbJQtbpIIPKNrL8Z3j9
TtLNabuaQahanEk69LcqSRU5giDvpn4L7iqWqAaDtmxFSOaN/+Iyo/Oa370Q7mKR
uLkxfEwVJXs1CylBHDrqHvgxKpxI5G4V9prYr8RGU0NhDPpwFLaIq8kstJ+7zPQv
ZX4BvBoKGfzM1CrCAsk+15HZwx97Wdu8uWqkHg9OSkgx9eBcXp9CTFBdnjkINcyJ
gS2+LVPS0fOAUCZsVglPryRmeW8mjc9xxdnAcWtcQ50xdNId3OPEx7kMww/zr94P
GSuirU6sF30G6BDGkUl8Jyp6ISQlWsPXeoIIE0DbdCOhAjEBgF4uEdqLrkaI5RMt
WKqOmEizGhJXD0w/uazMCcbyWrP0BotFHIK+zR1FI/Asz8EdJgU++OAYK7PlphS+
rGBXwcE3kf8Skd3wemMsUe+7G5ix/HNIZn0s7279BZVzyvNCAbVOGcFQ0zUTbpOK
Fn2mxE42n6CiuGYV2H1Bgj/BAmzb5zDV491DJck4iUAj00jOP2aMH7ft+UbMqxT/
gps+sM62gfF5MhAEcvDvHdg4tAvT6MXAg0oXZrooGBMSqUxqzz9Gz511ufnIejoT
AOMcfclQ46kGwdupBQhRDCVTjBnm1bM6N6pABelTwhITFgThvyb9mGYvP85ffa0x
69tdyLBDkRl8N1varKtLZ3dY6gQfK9frJQoZiobej41RAkTWGn5c53PNfBtWzR41
8hTS5k6/+fbrRMb+P4RLITe7dP7RSqsM6QXjqAN8C87/SokjyD1af4XB6go7OzJI
McZzcsytFwYxJ008h2UbVUjsCJ1Vre7lvWY3zWNDLO0wmyBl70o3CtVLrnuIVW74
ERLc2ftbPJV1HAGc+6ozNG4D+jfJwaTdvw/BplsVD1Xdd5HOuCSU+9xkDhABeKpz
jyHCDKlZXL3y0odQlgLLJv/0NxJJg/p6DUZVFOFWKdTK36ELxKE7DiDQq7keXuUp
o3It7sJBFHdL2QXvvNRzoysp1UAUCRsS1D/TcUBxzZSVEEbXxOH/swF7N5tmvbjT
eS35bNbJ7P/fLXwtAhvC8bSp6p4LNkjUwIK9lMl/maapMhM7UL8qdk1AY4MWJ9Em
ztHzjD+gYBMrgqJCiQ21RHYtqTs7nX5nCg76FmmzvisPlY4KEQE9LA4L686Y7ZFI
1LAeihJeFAg5DHtbxplEkBH02T1FQv347uybHgberssxoKXzueW5FWCFb8YU5X74
OH42ZVbKAvXRdWC4nEiBC82AvkUdMxU2erzyDtqJo8bRlSQXPNvhkGeRcwyGQV0I
WuWABNRb4NyXRLIwVm3LTJDKn/PRCi+yQJtwS3uXBLCBriooZu+ZzgUI11x3sCjX
vKmOV8/jN08/xImw5dGJmd/TNpxXisDqr9gNXeGiliY5c+6OwEqN/CitmemMc/GD
+/PQQgN2o9JlPIHa2gupaVPlSucj4tCLNo7RdKgNHcRM4cpy4OiXiyUTegYBGXvU
NozTFZ/jJcBjrDv7P202PiZB7vpbccQGR1xzsc8L1Ej/Le19Z3+lYRmy7nYiskVJ
0BazcnvZc54Sms3Y0m2N9OyAacNYVOI9ECNAmlLsaWpOosXXWflHhho51DJXxPx0
Qi7HfWsnDMuy2pgnSOasfzdlMUc2nYlUYSbQADZdB67Qb6SCjuW8bIvBDrNdBJeK
jGb5iEJzX3nyhZaG7EBT5K3fg5FRbUKfM/iYw+B3QMsarlhaDxsPcYgag97EZmSa
pczrQ+td8mCIdxYscnS+/HgwgrIt+fZpFc1lNFtHjoVO3aeMHNIkeD6MfUI9v2EC
ZAkLC9M1b3QVQKGDCi7ZQanVni4c1sU+6pdFE+iGXaIR2AlIoztzB/pEdLI8FsHl
Wehd+Y9p4NxpOPlV3cns1DvaYLpadeGZq7bNWGSb1WufGzCEqV40duz940HZyN9U
UsxV26jlau7kGupC1srBnaoJSs796wvSQZ76wQ05Xjqjvm/ujSgSpczYcsbuP3hb
IXqCHrdTXy0AR0ZKCVQDxweYHvNqCYgoVA1gLciWOe/h0jtgonbwysL+xHMOCQlq
olS0bwsTcl7s0chI7aF6lhfWRh2GiDx4l5gF3onhEp5tmU08gP3ulspjcuazxwjv
NjHXeT44ArDV6s8DXY2BZZiMNXNaelhf06tFE9khI2PWbRiOczZ4w7jCYC3rfZG8
ycptXh7ehC/5KATomCX7z0OIQDRV4FEoRCoGozL9mXA4C2ni7Qz5cnFjS9V0v265
KGOlqdpPbcX8O+ivEsC7ie3jrQeH6HVQSdvCliacuYPvlgDpVUNzZobI+3xSF0ue
BvcdYzcFDmQvbiOWWBvyL2nSptm1Y8kjs85w0zEFmaem1bwVkfxVe59puNNaawTp
Pt2ggRON2jMuM5Abb8sSUJ9PNt/iB1nOGO6JKLXlsDApfdyDXoP4qSkW+DWFFOE3
UACcj5iYmFkV4oEZRS7o22XoIcmCjIu3kfh3tUC6yekOkpQ4HdcAEFZ5od5dPN/z
p0lpcFA1FBZM1CzZdHZeht6fiRUUmLhTitLKDU3teu3Ubrab7re1fL4tjAiGHZUl
8RCN+mzn2kSx+XMg84iGllkg+OVTc6REvyWDTk7qm/XhwMTl+lEkdZ5OZCOGl47Z
0SMkbhN5lz/zo8PJL8mpf5pizNDsZuAqKspgbIQtCsZOksUM3LLLR9/8ZW5irkZd
f9ZD30D6C9y9KiAyFzmhXmImkkJhtBGheJM72E1PvYVazXDP3CInWuGFBr0SowEh
HymvWYn7ZXFc/IfgzH+hVpo5vQ7Vj8vDKPxxXyA7bDM9MYcQgwBVhlucE9M++wyY
deQkU/2l8EHYyWZOk9F/A/ez5eiiOkqIXwOMeIBBRY4YgyRanyTxt2cHUcMuYTpG
98Igi782nPJJ3C7SsypUo9+iu5kEgoPUfJN7rAFrWNzAAEt++2HgYUm0JZSNUyul
lIB5E/FUVveJ/45MpJQBdphg71eQABs516NLCgHcLm+XnWFpl9qt/g1iKPhzpY7P
/QmqJwWFLZ8vkie0Rr4S9IG+wCW8c0yUxcSwIvpGoGL7ng0HAo9U30UFyviOPreS
87tfwEZgvLv57GxYEbBsACKFxaSbD0T7oQQFxI9WCRxLhg1QTwK1HsyL6ezFnfGo
rzzvVwGTuewQAlbHHMHOUcoOBHLPQgf3CfrAdzYZ7RG4JViT4/xso/vnbs9rJp/O
BClWkgMGBVo4olJ/Ycj0nPVTpmKEFv+CoQSJdOskTAHEFyI6m3n4IMoRFN3ZInsR
T9paJ+9PQWVq4DUy/ZnEZdVyNF/zC/0bg4NJeFPrHH9myF78EDNni7MxP0shHMo3
QxN2crgf46284xqiJcN5OttP267i55FZxD8AvDJZGq5ORtnOVVP1RLHyQRlO9B9S
xBK39HUtPs7GfVkfvNQQVr2J1yBGFfxk1Yap9Iy1vBTnEgowzY86wyV45xR75aAt
T7Fk+97ENWkv57KPmfBk8XOFkawjxcxlSe3zfQyeFkuwH8HynJOe+P1Kvz/m8e9n
fZqccMOFHVd2f2Wp+1A50Zk3J6PJ81BFfaWQFweCV6G4hhqYgxIIrunHTbYQLdHT
/Vr0Q/6eAVe59IeZDybmZdMMceKGeOu6nWRbVmz/LWsR1HFNqHCUkVp/xxgHmzue
h9s2O+m25LknXaRduhGzZA+XvYOo8jO68bJomzBmpS154HWf4yzwDw0A0LrR+oqd
76jfKeo2DkJAUf9gGbpRscniWDNh1pwvke0h3AHJR1O7mJz5hHKYu9Ok9tBWJ0AJ
cYOY4dnNnIs08mHZVlmdPhgc1aTQfnoJED6rIhGVReCbFOl4ri6TgOsVJwYG6h6t
26bx+5Kd/blhniB6lu68YYN0jTacjsPIgzQqgJRIIGdzwGolbzuoa4Xut3ikQ2Xl
IBvlebn9v4Fh4EEmhGG46W2Ecx1aDwfH58aSVCusKGqqZQoBl/4dvg6KH4zyGV0n
BbaEc23Tn53PCaFb5zxbyFdOwCb3SR0Chysm12+YLbNZOxmOK8vx3IOXMdcDForg
5WXExq94KZD47PjzfkumIVcKigkx6mKqBX7zzGwQkP7w3Ia3w5UMkRC7u4+7qXJL
+aMakR5pArmRTiA1YAT0Hu+bPcbc1Vp/sIMRtyPgDmqMzv/spsdqe+j9Hc64nQaj
8FoSntUM0B8UwNFAUSTd+5W9tMKig9WGX0zCsDuWEn4sL6kdXBKUTZgfYB+aYjQh
tUfGYjNa2z7sCu2K3hcgg/IkE9646FT5Ix2Tmxxj75bqBUsX0RnKxh4F2SSV1W/B
qCTlKQ5O+T15peV1lKEPu8/WNiAXviwwhHnD5BmH5w9so7KAeqYABJU0zPflrExi
rPc2LXGKEJJ7odPANTjF8mebvVn1NO0D6XnA6hjw1dEr32Z5zwu3l5XuDtzljQqG
RTNAueFIhOHEnLLHV/urbO10cLwYHgBz7AZXCK+4lO8mxpMmnJQ5Kg1bLa/AObB3
mpwRCs8wS/mayslU6JBtLCarDLjzIDFdr/TZjLDaVxVRX8rFI6eNY2l85b9tqGOR
tbc+iLw2zHnPL+/b0XuuMN8lNQUDzkR1k1DzLVgKuG9U/Snz7Y/TuznNIUgpb8xy
jfFsIIrMl2HVD8I6nMHfr5MFFWHvkKdon3GMShe5/S14SHEQe1jDc16Y6Fbia6xY
8pwgbxYYusrhjN7gnpYIKdd67sMzp5CuDhv3ndUng2SkL4WSzCg3avjZe+d/15sp
4El5sqiXowdiULC6b3vUdGECYq3/sNBEh1bDWI2NzkhHZSvDzBpIY+S/BJG25HSq
LJ6TSSPzu+pEiw5qUWVEyCoOo4b3UjSlb9a2tn0I2lGnKaiAsSoRjFsYyg9Bhzxg
IUOW784mxgn8KcMQ/1/HxaQIbGIkKj7JsajwlvYh9kI50179pOtAZ/xHlElPKiOy
NrbH4GHnrxctrCjpC6iTU9yq7WHjfOTfanteK8f8yuN5Ydy+cB4n/nCz3M5yvS+r
Fco6r7k0k6IgZ+XeFMzjnXuw9pabZeM3UsIyJRGqsdYp207N/jZmX+ApE/Ruk1yE
8UFEdB6cR6olgdveaWFzDYLBEsH1tSvo1VMWB1bQkDfjA5mvg5RMMFr/LHwGr1Gr
AoJ1GKrg4bTid0DS5G///9MBIUM4A/AOHHqqDym9zh6Fdr3JJttfwiXeFU5w4mUt
DIDQ2r6tD0IulifHZ/tY/K6I+AxIIgQp2Q26dnis7gPKt9kc5o/gfqYvvefeC/eC
2eHEglOciT08kKAUu7AogBb3yj4j8rcyk0XBjTSWVIQrxlHd8cFIpCo4vstHgcE4
fBZ4rnHdPFAnuuNlb72wDI171WWUEvYxwF4LqtU7FNUoC6VN6EMg2t0I28wgz/HV
4mp1t4BKbuiOWNGu8Q143QJib6rdSNOGLv98gZpFxw8W6bfVw+8dRotGZlOfSWat
SmOqX6g9Spp8OlVJlp0A/+tlhPaU3irNgXBn/zJxfVLtA69R3mlxUPP2meALqfce
X2RNAXTGL7dAZPjnFexjGPLbdfFLXNw0MM4obdFzqva6ud1UlZzyPoOaTG2wvs0p
UJCLtx2RVx0KEJW+0j9Qx3NcDqyS/SwCM+Z11fKlv+jYRoM1LFwdpIpVlbPrmvvT
5rtFqt7S9ISi6i84ZPhhZ01mCJ9XbM2b6mxzwdkFB8wdosi1ZKoPuP1jEpsd5EiE
QzoUzHSy3wTFpzUAXkieYALWrQOzCGfkQfbJ+7iFtHb/rkiwi1AW7+gBfH8JIWXV
xiDzFl49t/fOZhdPbiSBoBeloRcVUgfbbU8nv9l7/50cDFRupYkKg7wyD++8QFRE
UDDnAWaKY9lBrPVGqr4lHD6F9zceJ/S2Nmx+gWCTccwBp4tVz9ErPmmCema++vFM
AH+wcKKWMOqMHvMjZlWWMu1+5M5LaFa6OQyL7u0NecJLxlz6zdEU+BMraRR9t0w6
O0Kc+qNpbbY+f1NdODx88pNgiQRKwdZXtmVE/JHdhOlWYyJ/QE/6ty5iIPNyCwgC
EZhYdUO+Gl5DgAj1TUEhnAb8wbdRprUzuAxS2RCjFpaeKi665ONFzS5anWf9dzUf
wjY8IHTz6HCGlHfGnGa/AULX6518TDbvM2ONNR6ZJbAmFJiwHSQSzTQwv2DhuH3a
Sv46+U52K0jaFMWr277LAblu8leS7TBnktIcUJgAPd76tRQUFAAaAsA8rYnYeHe0
8bo8So6J3xNXXr3bQuM/uy8EFvokMXcCYkKKhHmVdCIdzKizGkXbhr5znJIU7m+1
ifsFe+v1h+kx3naoZb5M1XM9uHXoQw5px8FvanAYFE3z3HLPvJ2OpuRZnaHt5vcz
cmcAPzvaPSWjY9IKyJ0QZNMwXVeNQhPiH4Gk4RRrMhCgnPLq10kYjs4NqtjNXQNf
od+GnxjG4kSPT4pIUt4LXFK60IacCVtxhjr5jXIu1BoKc4KYRYveactt9TD+AhXE
TLMWzyVvZMoCUHbkzHYrQSWRuESNOs7KJVIwq5SADzR7xICeBFqS+uBvab8JU/mW
ALnMtkMBkS1qHkbjbbdg8GsAJ2LCzSkxINbcLYm5F5p3Zn35o6wrE5yw4PgATW31
hBCxBq6VH7e/L9wdtGs5atQ9TW988fK4QC/4dfOAJaCwJQYQ6PF9dHwgKERTJsqG
HBMgRyRvRJCFRX2tvB3VAtEvR6l0Pksd2H89cfy+w4B7vo+JdNXKpetM59JfLczc
budOPOgxnX3/47X1WJkc3bJiHD2O++X9/LycdCmmliazqkzPk2XDTbBXSVjtlYcx
fL6DZxoa69mM2ZR3uHnLOhfOdGG6bXUYk2a+Y9pMqQfJFoSQsdLB/g9ALbShUZh8
+4Mwui0JLmJtkEIUrRpkDznYDz3KG+8j7hKlp42htkzXF7wwszd84Z1avU5dT2Hw
M5f6PJEduKH7hGVBQw5fRctn481go6geeT4wJugxcggX0XptSjTAKUEeo8PWOhry
njeUZFV0KoTNEYqGVeTzNNtr1JQ+Vgfj//nY/Ow3IFnLVwdXVy3pePDFaH6iXfo/
GULqXluwLb/84FYzfTpRmY85gWY1yz38QltMCCmjHLfg9gcx3Z9NizEdyYoftVD7
ReiuIfAmzZD9OiVn5f+bAt28bx1nF8R29ztm0KbCH1rGEtgWpXUdgCC3bDHWINRD
wWKy988BAOQVIDMVTEckwJa2pcVtvioxUraAEiTQRsO+WU7V7xDyu9IWEkIfL3vN
7EuTFa6DY3xcuV2/iGDF/TOFeWRmcUdlJVHLeAENZZKZpyJYmQ/4buOPbMvssu1h
aInl3R082VfPIAyuowX6wIu2JvKFr6d7/kNBvEZ13MEOtcQRhodCkJe8whOEoogI
Z/qZ5CfYT1n+VGxKykDPiaSwI5UEkofSUCA/UPrQS52wNYTQtaXSFpg3yhqKAgWy
j2fSVbxsYamv5kAdphOlB/t8+8eXVDFgMlXvUYxyNbiPYtxfl4DOm5l5OZyp7MPd
AO5nAzGkXaH34vuBWlYMf982Vtiv5sC4DaChzGLJPgC90kq9m8dviFEwn9c9QXfn
qzWasvuOVLKifO2Y1bWXHoqQ7pGJ6iPeAsVQJHpScce+J2wuhq34X8kxqHQJTVef
QZiHKr6ar4fcAElGH9oKl/Hu2DlKBsyX3QxwPDVU5QSpSXFuYOnpl4aW9hUH6yp6
OxXuhW3hYhn54lNF34YkGsbIKJntQAG79NCzQQFH62spELsWxh38Oa/UgpZzzZYM
SqjgqFDkNViypKbpI5rm2n3XVHECEfhqlJQ//23CbXKQFz+SAgP6A2koJiiy8shU
lj7Km7D8UUB+HwXdqEvShw4mYZTgDveBB4jH7+3WmUhp6Zu9EIfabj91Zpq60Qdl
5iMnPEAezvqm6Xf2Ehh+yoqE/qXQJeeGG03uZPJKQVJVfI01HoWOd9gpOKtoWVui
QwT7BSF/doTsl03lmajVvmZfn/Rml8dfkU0fCVijLiSX6hUZ7xd0+taJHR8Hxtjs
8+YbkfIGFXFoOSiuywlvjor0PH5wu5soZkkqvxeMoB9QPX/Z7iSL1vWmPljesfCV
BRJrdXE9H3LFUJwHZPlBBeL6iT6DQx3RFHRRSOfXhDmv97Nge8kfOqGxS9JHK/Xp
ggzDi1v8kRjzcehbWpQenC+Yp0CGPd/Sctkcuy9UVoM/elqgJBOW4O4XdHwXjTeH
p8nABoNvQMbQR7eOtaOwF0nJaMXJIWQCQDJRwMHwnIjrWV87XrtihrIxZYLGS5Ac
cZV11ZMD4MJn34GmTVO0TX39kvYts1qPw37Sw2nuV6kDKlv4H9eg9LkX/aOBSnaf
zTjJoYrktvXAiN9XJ8WHn0k5f1I/BmvBuxthvJ/E9QCOndMiyXrs3Y5PIZf8ETqf
si3ABueisiDTh4X/Uw713ZVy3weSFtnnuC+rWRU+QS6BpQbd0xGp+TuLEPnwGOFr
i+dApn7WvKaq1Q5A9LJ3OGhv8kFT/BZZucy6jvvRCxhtjcFTUX9U3IMrNv0j3CEE
omH496FIge3TeOyUkSRjFCCsAzEe4hBIDQ87NwbyT6Ij9t4QYZ1phOqwlAXNC16a
puUkFV7/UC2pU1XfWRjO+DEmZfUV2ZhcjgbH+yn2W2zRIWhadqQxm8lSYHZLCclU
J4eoyHet2Cn9Y4SPGsUPBVOx1t4CMILkunxgW1eiSosGbR95t35vQcyhb6DytXth
ssWcEJOM2kqSbO9/anLWvY4PeJl9SVCDta4Fqbzt8IuXn7rqXFhRKUKj3/SDkFrk
TKW7+WJS/N6kJYtEo4kFikMBA987zK+SmYcZXz8kR3Pt0jCwQC0RMo6blHluT3mH
kvmjVqw5rccxG4ZIp3CXTvh5fHE/O8AIxWdiIi6BFDTlOuN7yIQsQLfNgIRFtbC3
5HS07tRd/FScjg1jS7lWX9KWE78gzRZD2AfbQHR61y3ck4R/mo0URXz2vnSgBb7J
zUtPEbW3oWiv33RbKtqpjRQyBnvSVDA+6+mRPxgYFyS99MJWSVPDf+JT0HY5tax4
FWmHFFGd1ic9y/7rfxughVI0WyGd9VateB1m3yB5Yr/xmhdIax6udi+7ciGEwX12
IslwPkqHwixyeRLbqBULA67VTB3ufDs+2dZs5scyRyPq7TXfbVdsD/9QA6RFepB3
FlNSNQX1dWY+HWsmo83TCFCo6ydKu60+v/DrHYqiPyEJgG0VbOcAVy7bdJc4Ug0S
c7LqTfhgNOjhz0O8QH4oqCnd5B+xvgyzFAfohZy5sl2bvXnTO/wSRUjD0TQ65uAv
MkTTwOZG/6jDYXRRQVx6xw+9aUaASrfpER2b3Q7kR7lkT7R9n2xCVkaR7/rPxTQ/
HXeeJWjYccSm7er1+Tmgrb33LZBlzQv5Ehi5LXRdO1nDKnn+UfoT8rz8OcWPz63R
lB0EOy/IYTqjX6liIoA8hAJ3asIWTH72i49RV7809ynNmKYBydTZ4GykO85KiQt9
bf5q4VXj40ceWG+qNW4gsepOARasdxkcTNmKtC0HQLLtwz2TuxVQqDff3B6oyI7R
BYYUKAmydlfog02Xz1NrXOZc8Uh7hUnvtYPykr59nDxgX+3CBDRiPpdA+de5Pxg1
ToOT96L3hdI0VXDkl1dI9UXGBYGF9HkAOcf0550TtIsS5wYSbKDDFg9oHeu+pmUp
LlixOPC2Tvp54HJcHxLLbP7s7iB/ztFBw2D1kDHWek1+OXtNlS/SnhinGhUOV+YJ
U9V3gRCFU/oevfo4ZBtsp3fIdaXPZZC8b6zAcBJf+Vv5Tv6o+zqF25B4Jog8UUCx
4605RlvSIlZD4eJg7/FYMNUstvwfVp1JJWZ9fO7GQ9CtpWs+ah+hCxznsoJyGDiY
fgIlCek6t1H+GxWee9IbcT0rNv7HI18rSL52MFO0J6LdR3hM0fHwBogQeu4wpFUU
goNpBSJiXLgq7TbSTQCH5pht5Pa+SxfbQ+K6usDrGsaG210nUinX7DlbuaPauIoE
o5h9YYe+72hdVUCSzObF0/lIrRiTdRrXk0/M+XwKCmkzb5qFCFjGhknWFfEJlhgo
h45b6BbIwi3Mnh4HiKZr8zzRvWoT8QngLFI4nPlnzuN+YNTYCLTyB0TQqnGq/MAB
G4OF8WikszAoe37S/ijDAMkZ2DkeJqqsaU/lNjxIJ3+GnvqL7hHHEsIF2dPwk3Qp
DcVUG0X1ujayLX9osZabTzEFY1PLqqwEmUp9MdQMG/Ciz/kyD0jMsRgIdU/ghBxi
D0rNNMJHpnEMc+h7mBNS6+5tyU3g47pyzLoqEMNoko4l3YKHw9ihs8b/uoK9ODS0
HKSxnXoztXRXSenaG23SpR6lZl4PhNb6SYRXM9K2mzFAZqYuw9SA18C3Q7OSKonl
1EqwkENrk2lNcIDloc9qyx0z1G8voJ2RUqgbzIc6ticTk+czIhWEL/4qGDo/jtLb
TxDTLSFyYDwOKRlz3xe3IvEwHNQqaHfq6jvyusK6WYI87vwMJUUZqAI0ORm+P/7P
9rM7Wol4Rk8fDR9qgG7id2UEmauMcHu0ZHVoNwXoa/AQ0oWx2Rzok9grTkKLWIMl
IeIkjemWDDCZF7Oo73v017uFSjqVGrmCpS8uKAATr6mJ4WRGbp2dZ3Uke264OR4E
/P2VlV/15BiGbc80UYATwqFntBsoYGjZHlvIvlRTgCLwXbMf0elQ7hDhT39+PwnZ
BUr+aEwlO+s2ViZO0tPq4FF6g0qf8pYMStv/vXPdwZ8MP1JiMGj98CpxQ+gFVRPk
Og4vjDD7AzLqabohrxSfQqwGp1GB8q6ASP12Ja2JfVwwvz0SOe6gZ3llCCp4hMFI
7epCFkgxpUguP5VWKO+sJ/iYAYIKKAEy9lXzFePW7b+M3OcjypUF/lyWy7E+KFct
sttV67bVptdInSJL1Z9hR62ejBY112VTeIuMXe6EzNYugxSSa3/obXGCJF4cY9iM
XeMlW/5pIBF4DU+owkA5zFUPU4XxBiBXFDK0+/flSJTwpMLUMbeXG9XcX+J1uOYF
EnKNZ0AsP++ARAQ1wJd9B7nk0a/vPvF7VQxZhqtGTKPrO/5FzDeupSCM/CmabC//
nW7icdBtiAOkiWJ/ioH1blcBxW+RRFu650oSa9YHFCrNODxnGndg6SJuaYfEzcKU
9euwNXCt0WKBQaRhqdbW+W4zMcbTQSeiITCpadWo4YvtOAGFWPzZ+QMDqeekhA0S
fKvbpc2aj3WvzljzRqRjVax9Ec+JDiUhHErgC2xPd2aWClNEBRblUalXwmwjI8mQ
oWAYwQxGQyGhTukixGP/6/otRJWahxoXkW8ej2e89epDzQSOBjpWrdmAOQp7QEMI
kdcO/9Kz7xQ9UIvzRX3O5oT49GwkUr0N7Li6EOXh1RTr3UWEl0oxAgKrVkwS0W5L
ltaPMJFoh6RynriYRLGI2J6iAEEYxJUxAhfQ9Kc1GBopdhMSmdvVxh+crmyw773/
7Xy613nDYranu12mmcYaNf+9d0uXQ4a+WQEvj6C1/9pLRNAA8dRSfHLK+VCbOspA
VNiWijn09BO0VBu+9gc8QYsHB555XqZgG7spdCBH1phVGzuT68uZPt1Ck/WRm7Ma
bi8EyWuelN4N0AtyjgY2MUIm51YLubscoiYtGkO8GjuUAalN2LX21yXwCIQzY9UY
1pyrD6mhodQuq20LN5cvfc1eNClH/1/DN08iK0sSI9I/QD7hu9JOD/YzM7Qkgrzz
OcMZeVTH5clsdD34FfrK5CfeZgH/3OCD7Tb8WnsHSFaF+wTERDwdanfYP11OK0BH
vPRhymH4VLOO08fVewNnuUCZRiknbvAKpefciIc3rvZkr0POAmDQ4I2W+yJZG3ML
l6inrCcBcXyvb9ky8u8aA39Q/UCO8U79NpjbnevzCB2YhQfrO/QrPl6AtZr9xnDm
dqyBaKi4Adj6J9eIXPN+UPCWBSdJx2Cr1Q4VqVCncvvgylsdnBVefVWXDRdxuAkH
FYG6vNzjHHyMhqubPI6JnM74d1lGydYgBC47zaiJZxZ2hhXZbQlP4DNw2utfbK1J
vDgeDQQSVMM5EyhrB7Vb5O9ZDjYBGLMbs/iQ5NDp1/ZyOCmozFJA9+UmmbNAIXin
pO+GrGNjwtdCIBiKkqBMayWSGOVYZtJZi65rVsdnQNSufF+esc8//JWmjfSBQM3O
qw9bejfHsY2BCVG9OFLXHeyhDVky3NErhN+nU+5z2tsnSO1RhQRF7vAcS0zTVXUn
bMSIUxAIO/UerAZffFvu3RBa+w23PrCSyKrD11cSElVVfZQefkekczWUYWbwRgaf
S4qq9g7kGrjCv0Ux7dkOVTdEVQ9O/fjNT940RlKuDRwdF2cYvdj1BICfhniBogu8
mqZlPDXwSzRjFsz+yNmHL6jtTe3OSHXRfZcjPsVanDEymIG664Zl36U/pqnBzetX
C5BP4hL+UwDeprPtk4GhFVP9sRz/VjO0M9UUWqvrlwmCOx0PfqqKRGjl/S9tIt+N
DzzWuLwt4pVYbs99QiyZzpw6aUDfJClPiDvafco4EG3mDNUiIAXuwcLrHDV+GUTw
hW2iZo46uDFcWd+BSpBT8iL0QqspSJtwWZ5FBjXa3X2ho/h3Ew2HNCQ6j6Y9Y78q
K/pPHTICYscDe7sKtGzzXRYbJFgY4eUFujdKq7zb76gcMoQpYxF7wvfHqjTEnqyk
E32y7SpVf8UHOZzZu5l63NGvDl1TVoCpmeedhy2H1E1DzEfIPP9+shT0VaNPrXJR
avveZiIW3OzeSkQWJLC26NJZkuTKb8ZUKS+E8VJ/P782S9i8p2VsFWLexCFAtM0J
bSCd9g1iSWE8mp4zJHiZmZlSFIPRId+2GBoOaK29YDKa0cWCdaFyyzblmCIC71Op
XEUeisMXs4xDtZVRtyHTlFpoQsduWxe45J+B9r6xmhq51dSNrSxx50Aw96kI3i0i
JsJia+Fezq8W5wFFmBCE8A3iLvmMDlms16PkwE75NcwjHdTcYdAOGA265UJK3KMC
NL8xIML/JfYlyFIEw7wbm1TOM9yCFcNzozn2a7cSnIO6Tkh9yr8H2t4mdBX9F+hh
obafYQ1Oosgix8UwAoXuaA3urnt0KCi1fXdL3Iy/T5Y55MMEbr8cUMtqlrCvAVoZ
Zi0DN0w/pzRBinFRgr1HFveu8sL7FHa71rVOqmBUOzWVxchmFpDbjb7pwV7vVaKB
3/6yNsSxk+UfCGQ2fZjDye9NhG8Y6Ys9ELWhDM2RLCfiowYrtIrvlhqHYvRvPYSv
LcskadDWRgplp6CmmT9EHYvodZ6R7uYpSQU+X+eOEoou6Pf3Q6/bEDrfgLs8fsWD
AiobtOu/5Ztieiqm0BioFwgcDeR2xox1NQK+IZghClgEB20eGf5vuJ2dxMctFLw6
afFwc/PgpVwXQXzDrBoG/TGuYPzW/JcAJ/DqhMNPVLNxoxyxe12607kfEGjQ+1Sl
QZlQMatB9HcS8C7BtiniXet0pl7GZC5KCzodi3e/wAbOfCqT5boAF7uxSV/hPU+W
wl48PFDHau5eIOuiCwsiXQ9g6F83gJqYRLtcuR3AZ2SR6fkPqIfGEhy4QyMXetBS
iHPoLOA5/SxewcQuZ8slzqRIuVFJ7aLq3YEQ6vpxBi+J18R7pcQ4UmN/k62/KqBL
fS6NYOkfNBVRAch7CBQjZbBFasmR/NrOy1G533ootcNgSKS/rjbZm+1Vn4Y+l5nt
XCHdag2KoiSUtzWBW3YbnUIYP6NOvaHwxdzfG3qOI+UqMvUN9jo7TxPkm640vxAc
Qa3SuF8rjxMeCIIJ0zsIXYNZ0ehwIPfHIbojGhwmne2JpAXcp/SRBSIIue63Mvu+
v44fJZTXgfJaRxAOtAV1mlqZdy0JwFNKr24t0TOmsinxxmpjRjBsoWih0eFvVba0
qVbVyKWkATcjJ0pNCSm4JMVMuOlTb8Pj6RiwprmfBvGvAAFsnjwzWNS8GVZ2OAam
MezgkgT2rocsf826R4f9SegzfhRUBaI4Vot10iRvpqr56R9MZPoH364I7uF8jw4Q
zqpBCBasRIj80grS+czbi5J/HJJDhU7nKGk5eF9Pd75HxN9brGA0TGV1u9rXGLsq
bOu9CvWuRciCk+dbGD7NdP3vRi1H4705SDJnn2G4hhufOBmVfGtmUurjsDmeHwzT
0w6pX0qqXc2bUQM0QL6Z95AFq317uWxBrUUt5/PVVszgLnM/YxgXYP1JM3iPxHwG
mZc4/PoYl+ffztCbgcner1oxZL9rYc11Os/dGVnHd6yD2ub1NL16IPtaUCtowGvv
MJcvKHYDhlvr2gTzo/iB0cq1g+0JS7HibfphRM0z5+0eOOn3t1+BYmUxZZ9irRnj
KReQKkX0THZ5QlJHMZAAIfHbJVuAS1tu1eT+rsK529/sZ/eBbf8QWOFYIj/jsb7R
ovYf99WkW4hcYeo94dp1eVrDLniL7E6xW0Zw6/2hgubBsXBXEkC/kolg8x5ayJN+
XiRjFn+5w+LZ+Jdxhqs/eP/JudLj+KqjKgK6CcJh5sgZZIO4MJWo9xpvzCL/Nj+8
G2vQUIaiOnJ/XmdMWXt6eF+Hw2eaIT8b/3A21pwPHassUVXGezG9tDIo2kf6dHus
w6XM8DfjuipGK0tgdxv0zsl9XqJk8v4PZbdTDtRDFRaUjej2cF3gHlcPhpGcpedt
Pcm2IDpfzDzFwkzqGkdP3wRSr8hstqoPu5fyl8+eBMwgr1EYk1ouWIEXg0j4wRBe
EzUSGQwu6Ivc5m/W3vSA+45W7TdTMM0fZUnV//8DR2+FE/V5/x/LZQLBbXU8i3nn
lglNHm+XgzbRKPpFGG3Jh2njOWq+wmuSeka0nKkOMv5i8Z6dbXQbFCMklhe7j/vK
TWNBGuHSM/Xc99EamqNU4pszkRcvtAlCLfJE0W47J3qJn4+sHjjyEb8F3ts3zTCh
5tg7ZHnMHK4EFGHCTgyaPuT4SeHsn3NLavQVUvGiMemHKXXYNgpzPzAe1kTmzVYo
tbQc3fjZkoOqYeD1NNOUDAuJWe74/zSMQ1mhL8WXaTBucLDKe5DIniuexUIc+Qfp
KXyxZt39/zhcze7eA2lZfcCHq0biDZ9OOCqWzR7jYPy8yqyE4ylrVUtmMMfljVn9
ofmd+i7VWN9v3nWIaXdIjtXr1i1lVUrTVAMqBmoAmRFRolzn1JxjbHfragN29zoS
0/G8MWiir+miLUNZeONy0U4TLmXOnsaiH4TFEKyVn6rfd1gRo23GAKIe6+G/hlnS
0QC3sEpVFvyZKitu6XUWvpAAUT5RL8H+N5+FP5UYB03iPCV2pWve82soto8q78qT
0QnW1gq/d8UmWCLw6XHGbofKuoRB4Es+EztASJfSQ47UDIHv+D3m9bh32ImRC5KV
zDM2Nj6IUuYflQXbTdJu3TTiXgtSmxStitiAtTZjKmey66H2Hq3+1mH+h0k9xj3L
EuNO/U8IYBCTfYwuU35wWRyNvCrY6whHa5rV91Gs1Wf1TWIY9clft2qHZ/R9HAZm
82LrfWZdft8fuFOjw+HXCkDercH8mxLYva8TlBlNjbCDojc6x4YvroqdtKcxkkA0
Y0x4mB3XwzxqKYiLq5qtOt29xjqaXlFqZiS62ckPjDBrs5uQfjpWTRNDKwGEJs9X
Yo+S+HIYVQxCYU5wmXh/e4G3RSSeUkVpnKKXQhrZT7KZ4xzLV1u2qNdMiT/nTB6s
+4VVEMZkXEpsdCFP2lDFDYyICK8Hc87hvFZKPfpDVH57GzcNLy+YEnERW54bzr96
5Xg/mxRqSuwAdusU2yuwQprst8z10/gSToGmHJ5wOn2nNkU+0l9P5t50zmkNgIqy
9vXqqk8PsIyM6ObFk+jaFfqm6CmgMtSgrD5k9xpfproudj8b6VyJynqOhxrWiUeN
D0RAKlH0jqatEiOmf45GAnKK+zShU7Jlv9noDAf3A5EhCSBEBU7405A1ZPEzP5Uu
xmfIuKTQ6P0ubppLzGow81KuksKkzW2+qXoE+5OoNtC2jLgX0HwLTCnh36786G+8
PBMExYcPKf6FNJnRr0jT3kiTQKeIWqRTv1Q4RsBRDHjtKRt0cB20ObJXquB81K2x
uiSccRUaWb1+RvVc/LdJgAF53SIMyAQ5L13clhFnjfF65bQAfqG5ScMLaaxDSX90
Qip0w7A29dKH/zrHy830IEAOHt16vX0OMYaqN+Zdw2/L+7jGOtGd2znxxOEv9NSq
QaysAwqupJf8Iqyv98Diars72iQ+rmcEY4qMUPduofeP84aGjkugai68ulT2V0w9
DJHRScCXyJcxXiyiqxaZJC837VPOoo3CkE5LDWR1DrKpsCq+wp0su8uRS1mA17EP
5rEw5cMDMe9ACgTpmmw8pZ857vGtOsKu4JvjVMTzRVp+YBQrShleZFS0rfQVkY9x
xvIUwF7rvuqmfgi5K+wiixWufVbUQHnzphvgk2GpuFIMk1fLQvA8Fm5mbexVQlgv
00rVZOc/8a8N1OK8ueeVglBltZefoH5udJ0QQhlmIc8eMPlDqepljBFthhMDT56e
719TS7BLYBKA89oeDQ5L6qfhAyU26bD+PgONM1i4ZfeZ/6y27sW5nS9JJtquCMMW
KBX0Z777wpneEz7DA3xj0DphAxjqWHdbDloV5LqsDPlGLR2nFo5NHWiLX/lG3ymN
VIVDFG0c4T4IOfl4F6Evno/W5PPgtwBBt5/xcHwpeld3ChPGeXRMYA7IUmqW/qr/
Dct5JCypPhN61p5zeMwzIWIdRjQ6Ha8VnMi0H3T2DTEYmjD3GRiQRCad+LmF925u
mVoTHBgmht/yGVbhg4CuUxTJir0n8vh3b1KFxXCUubOdcwxq0xr2BcYJTia6UV/t
jP7CXfnZZLK14PMON6GZ2JeX4/z6ZcXICN0GvsYOPJbTRsU47L8uNtwm7+CNcoWG
2cFgftcnhvvJZDPV865fRXtU0y4ftSMYzuEPp5Z2JdYfqpwmS7ONHJcvKYFZ0fgi
TtCO4K4SM8wiC6E+V/Kr9CyYNw0+NWSHyGux5cnoCX6v5V9z7ktuaLecvmPz9A3U
blD8kHrnmYrB41HI3MrmJwrcy2v9C8HBmABSZv09QWOEar8GNzrmLMQpDSaf//ix
UjN4Qgy49q+vo6UgG5G52OHP4ws5NTRDtbRwWKnfVbfs4ivoyaCeHYPr9a7yld9i
OCwCvGuTgDklqR+3F8cokvp0WVXzZ3tTkTBPo2PAHrtdL3uaPOVKbIMP9Pezh90b
N8X/cBU2B6nBwY96KbEz+X3eI7mBEhcHao1oo7li0ADtci+U1fje0h9wLy0mYNmK
UrfHvKMXFS9FXdi1EjFdsa0PKHtlGxh9LfvgaPDLp8DHsbq1/n+9VPVcTtl1kQio
uiXV/nzBZnuaKSWtmwLVN3Snc/Ybz9HNmc9qYDOzwHy30kI+8FGj4o+FXKL4ernc
f7rAN+MhSZ3DDY9T4y5pP8wQaIW//B8YPZPRIVWjhyNCFPjlzI+SRkX29lXhmWdB
2BJ1ABV97K8kohqxyz9QkfwhDVu2tMKpxYOHyIf8hm+cU3Z3oUbaEhvWSDKkjz3h
8FB/AqWuSCHxPvEtwqwtmtNZiabd1+/C7rRjz2jg9mTc95XW0q13fkI6Pl1Vw0tG
+s08DBc0fkH4lPIk/h6ZGulK6a5dIhay2+DSisLayYJQATxZjvws33vR0ejJIzv8
2vm6XcWR6vDlQm/I4mkGno+DCmQMdP9FbtrioiAybyLLYoDh0Y1SphxIUHoAFiAC
3jUQHsubi6xxv+blAVcej9z9qOal986PHGnCVH+C7d8aPY2bjshcrnr97kyO+SyF
CiScH5VeQsaHt6N71WRkSqwB5fwpUjYf305H/BSlAyPun3ROer0Yog022mv91egW
QGeBi1IZgnHO4+PQsrnUvoz7UaSRNGKHdxUyHbPbLYSum7DCQ+uUeoBhIdK40b+d
slU3vnZAMTonzZJvdHniWa0lSYNY/CHqe06Sl3oVZxY4gaPW/GSFcCTnz14Q05kx
AtonfgMiNt5H3Aad/4Kbt1McEXcx9jl5wSiOttEsOO1UyX9W47JIKeGQLAYoX9jV
n9616P5Ko14Luj81J02EQJqu3xonM0zRdD0ZIfJ5qeDIdspJgIzzDScC1raYD5c5
JoZylbR/YhonSjIrQRCrdH8gY7UW/uAzZD6J7a/HGRBJ0wEPJYtOr81+NznAtjuE
bdrfsc+IwHiRIClbPej+BZZdpJK14sgc8zIkw/34HOMQnoBO3i+uG4jWXaQUnH0l
VPeHJV89Dj1GBXjMutPSW+qN0XJaWWZa5rd7HE+oQ2Yb0WThKTCqlDu/KvOAFEDb
Q62c3rk3qolBx+LqyLE3jKWQQqyqSJ1o8RocOOiJ1xhQDqzx7XKYt6eSS/6vhEqx
yVUlXpbRH0qfCbPf3pXnZRFXUAw7rvdDAZmNUldAX5jPfdlMhX2hctrhA5knmKzh
2SlRSggjmAbpfx3ZjDFkqq1fBnLRA+JJk/EgxXJ+syOAmIdCaGi7fOssPHflMYOU
EVwPk+3EwEj7lsv0XIlgSLs/pldl9jYftcgUgJ/dVEkBjCWt76fuKpeb7coG/g+R
PjBFNeSJqYrvxWorxO9MKuj1b+XP6DRl0y5gdY6wWSJHYMFXS8PWQaVofVejbdy0
cNjRmnWy623nt9SePaZMqLwxQ/FuPEW44BJ1p92ct56Aai9gTQ4Yo5lzqdau9cSB
PjUdF2sS8+oGJW87DaMdbGZ8kmshhb+U8nCqP7tc9diyP+2IxZqdmKaTZaE50fQu
46zQcOY6TkCwkQnhLvGf7G8453TKkZd4jspqJTcRJZnd59llc3E+AuagvNgI+48f
THugFlFfHe5f/30AOTe2W4yUHcVhP7fmI/7a+1Z06dwq7ZrDkVrFBxDW93xU64P3
xKRgP85+z5I7JnSA9tip8cvvEEhl4otJnQ8mmA8Ayn/w9vlR+Tpy9MuFfJJdoBXx
rUkbhYRfl+Whw+TfVA9k5S0c6IBXUarK7/xMZY8X1oB24H7nO1TH12TKnwffsQkb
JW/O7qN8ISdOqQL05wuu1ZIC6DE+HpXnJykR9igVT9VhAaFMBAIyG3xtVORqsLgm
KVoUrKnyJDE6VIu5mgvTeEkPigLfqiHF8HkfOvlLU+GJpQuGlbEsn+dDjKXjB6qY
8scQAGnqAco2g7A5yczaxwY6g0tWHt9nbOAgRnWosdJRtktvwmTzOae/ZzJ5F7hu
dQXEVnXjBhAY16WtgN3gSbXVxjq0pTuHVlE177IwwFkg1ue2/2SFVxIkT16TYV9Z
I3xqVWk0t/doacQKjIhLyLUCMuVT2SVLk2vT+e+CATDTApt5At0LKzsUonTcp3E9
6uyb8/q6Y5jIgkjL2IKfmHkmDl88U1cf5woRU61JWEjXb7yvxXmmQoz9OGcHqqE2
oXf3YPZ6eQEK8fkuNDlT1qnea0Q1hOod26u6yYwVg3+EUxjVyKhmgv7lRJcR5aVt
aJedCQ/g7c/IB+63mHKDq8ADb8/tiJvNSFqIUSLsNf02/ZldqLaJAXnxPOOl4EWW
IYB4xZImhR4wckWL0Xk4a3+dXklDMQ+EJlBquYLnzpTly7mYnumoUoQYd/BtIniA
T71MaH9f8s5lhKZPSx2AmhtxTayP6j3VXRd0t3TPBDkaJ2Fat9YDGC8xj0vfXSGp
DMD+I0zXcVoKuooeauiDdI8uQDDx2bxYeDMmQWIAL/EJXu+I/ZPpjPjqTKLDQPg4
Rx6E4muiab+Aak/qsJ/Lxt+2VISBMeYAJ2EPaDkFoeagsDR4CBzMJJUCr1ddtgV4
Ljxtt5wNhjIt02m8D8WZE/Bp1y5Q2smn2OAcjImflYgSvJFP11s+BluiVqf87btO
Uuc6pV9E1lOtSjsg0KN9eEEwXk8yJKdh0wzEnKgYwi2YWU1Hww0n7ldQEIeaHPIQ
EUv973noz1AeYN3WgkzWqjQuuVPPWqj/B5umQ0djuzJV7Zh77mDmofrVOJmRNwaZ
xqibSHLE4NcuXi9zlMexe3BZlb4p0Sx0Bh8LuldF0i6rUAhP3lvg5fF7UFvVc24C
9BNwkpxmGHgJn1+/MYrX/+UL51ti0nqNXD+OkaV24xwo4QILWqOiojGWKGtGVQMU
Dq4WulFyW8q3xmGWbXfY9+B00MeDI8cueuB6RGINLeWqgWqbjP7idqkUKDzStCLb
GQXf0jIE5bgBptqfSfN81f8kE/aLuF2J1/V/8Mp7xBnlajO/iWY5bd8rAIKZG1s5
GqX70BUjITpbraVEwejPOFgpjqKTYgPxd+Z8MLCsZHYmuLjwHa9jTWNYAgpFzI6b
OEIGpxLrLgBNRX+WN4+dqFmHfwF7mNHnAwNPrmnM0RAqfrk3S4k3y2D40d28ISJW
OzzKYxX+TtW62tmfq+9ru6+BjpPymteZCGu+3edXzIx34fVclDXwglB3GW3ezpQ2
Opnzz9Yk9OThlssGU6v12Aiy1uZIJ0BLXGw3JOWEnXOBaxrkN6v1ieV6+Hu+/hOk
e2xag3Q5gcYaaDbzMb6bM5EwLmXRzF1keqh/d6w4Qy4d2kkSD0MYrueYy5KxP/wy
UMpmHftWuJZas8Rrm0Sy3bkTg2qcy0XoB4B+9a8/krDxhL3/0Tr0U21GmhoxYHwz
S+IOjgtbrLPsUH6U+9j3H4ibKDxIRM5iNIVj75JIl7C0WElwKYibv8Nut05SF5fj
6iUuQSjFH/EovbpdRy0shh5wIWZlDwuTQngBqaXPKh6uXfSjtkD5B3ydgvXtwqBQ
6IeJxYDsZrzjVLJLAla+3wZ0GRhC4/8qSWXSENlzJ0GJgPzrKp5itqR/8rGb+m5P
W5poZxNqNXUDwaap+81nHjfiGVHfioqPFBMScBZPGGOFveTv4lgR+SjzjnAFOXtb
x+X+YIMCnxcAguUITZC3MTpF3BJngjj2bY3xlBft9eq8ij02IAlWuchkP4Dll/YR
X5NKSoLDU1OriTRfl0bwz6Uqm2IH6EuiS6yC4XWBPsznOfRYFYqr0MO+V49zrm0A
RJk4I3ilspe0wrQ4h28jSKXFyJpv4rKLRBoT8thsYJLus7LOwsgCY0EfoTTN+jEs
M9lcC/pZtleQkOYeudGy/nFq2QfGF+LHkGbAOVrE+GARJn8Q5Xyr3FBopapWoODj
kfi2I4NQw8BZaUEUeopV3f2/UvTHOZuxcvPDUnCcX5J8Qyw5tcPudpPUlzi76298
8CeYdNYJb4dhhVj/6K6A/AigwK+eBFpZxn6RwV2mNX/kN6S7z3Qcvw0Yek1ohzFq
7OenBbTKT3EC/4zuOIYcmT+FFFDuhI7rk1rK8iCgKSqpQvbvsxUP5wSI3jhrxxTS
qvI/8QYiLlGJImqjQHrYYldUrt2ilGQh4uFQgm9T1EPegFCkwZHUaenZoj7TVatP
OHMWS1gsVOesxXRWfDnQFiRvcsQ4KmkVEwlGemu6Q4zHRTEi0fOAv2Ayq21gkiD8
Ei9TwPATOpsMmcAWbofX2sTcBCtTCJx+hoChsn+in8S1Eu5sBbsTeJVum4SBrsZP
n8WKqIPcfAGU7zgzhuyU1RBnikklNgxdubVPcbv1rUTu70byZtW+7VUZyeHPYzVr
/OBhFPGB5+511sQ6weOXlntJ0Haz1/iiYOQLxfGDYoL5Ir8lg7YqytttynDiF+j2
C2XKuo/s8atdj3yuM6bTQSKJaaVL3033a4NAdh7THlO/D0XU+ce2tVoyxBIh5Ad+
qrfiVXQwdfW9YEMdJuyRK71iPLIoKI9LTqNL4+0h+uCzfPEtAcaTo6Qx8XIcFT5L
PVjIA2ft3p2SZK5KNDsyudSseoHt+9AOmk5TOIwmnKvTEtYKevPraBI1UEfSzeBi
rCEcGmShIw4ykku0j2YQfy62RZHGqZDNfOVbd6+/E+ci4zvMxs7mk8tTMIDLUiXp
v3w8rU5YlCARIqECRlTTZqK8wIzcuJ9Gp8fCpN28B7WS9eYSgY7EbZ7f7pvVCDi9
z6ISF6vykgPC0dASS+iag0gQiU5K2diq4WlxkU0CYfdEZsrnhxol0Tk/uv+V4a8G
Ip3IIkJ6TVVy1xzAHbFVBgHvVR0Q/xF+3uIhB0c+9hpFujIo13E1Uiqo2HK9f5aS
w0pUsntqpfkk5KEQPfmvJt9t3oDMQT6k8O6NwOkLboSl0u2r+CtHZPKGNmF0Eb9a
MQhHmIZrhi2TZmG+Tj/BVZcQagjm6ZTtCRMiQD2u2iy5AhPbeHDRUbUO20uKAhE9
UhpdSIjMHDuV3p3T2rF3/AkzLNbjcMeH4Q4JxICCt7aWzkJEt3fUMdgaQcBwbWJU
OQcbm3EaNliYqOuTYCypNMFoHI8Fs7xoNYRJg14aNzXgZMS99zfwaMIABTiDY45q
eLll9n4XHg3nM8PQRmMwpSWecTp3BJMsZRUcYdZZketDH7ehD86So3ST8i1rQ/xZ
bX/RlXoV4TDERYi6g7gCuI13xc5AVTud6rVl+kIXth8yXdyBbGd65OcPn4ZYDHEZ
VpxeZnDe/kSjFjIaSPG9iC5r4aDvcoUlN53doJsswY9yAozxc5Mb/K5DtOpXPUV1
LyoreFS01I8LXqHv5v8VZpkCBTkptZ+M3GWq+MngaCOtYfDmL2Q04uWGKE9p4IlV
Dc0YGTm5Nsm2IKgVbxWbn0TGtIP9PAzQSXiLbm+avIqSeyRkOxZXQxsCwR7b4Bpg
Yk71G97k4OqWN+2Q5qX4LwJvzjkCakd+RnAOxUUkKiWH/ICfXRelLxfle7d8arAi
OXO8aAZeFRgt+KkQO1F9paykhoekmUUMbXIDu34aoUf/nSgWLbR7r3ehciHeLRD4
pkqUWSL1MvtLRpswR3IdixEJgP579ggwnxMHbTtuXWlMox6g+6xqQ71VAXmqr6Z8
jAtABabJ1oVakBUgjhkGnIFD+zuDlADHa9Fain/31aQ4kz0DpMK1Jz8SBbxbI3+y
X6BrXyyWvn3tD0Ic9c38CXCiyRa0xonqkMziPHSWe6rAMcklwjw3NDDjJD6xV1Ct
BLOFWRvmh6WbGc378Ab1Wo9Y/Dd8JCHDa6RfNyhlLU1U8rPOetRf/FhmCW7V4Bdp
IrIq53BvPibxDNwMs1fE7pz1AR6CGkmcJbfrxgE7adQ93CNHNlgzl7kVtBqGmWNY
Mzbwe0NmQtfoM99+aaHcDsxzFnlcy1BFPQBNGf9lt/e13cpifwhWDhHJSWG28dU2
gZoGpUCxu1cZQcMpJwFsUzgXLnJHS9dArZilg7UuuX2T5Y9lZQhbpGBBZDU3gfyM
eXgvIxCVO5XAVX3Q6AfcI0/qbqlJ3nMfqX5gqqibnvCq9LFbXiahZK/LfKfn7AOF
ToNpJP/+03OTjiko/4PG8JGt843ashUqvXs5+ocTszZPc1eCy0n9lWTkqWM3bKyM
XaezQOeX9tvyonJyYvQ74HYeuv+53dNXfa+p9Krzz3vs3/Qq9TOLNDTRNxKsDLZe
l6+oFm0M9+iJMwrJ0lgVM0bpLI/ESG5nJtdCWBHF9RyZ4sg1rM6SRGIR4mZT1Wa0
i4XfB8OLuIPaXUSWjE0j3tTGvTjt+5elhQfjXpUZL8PbEQcIWTb34fHeQluMqwRl
NtGie839c2/w+3Sw5xZVx9ckYc3WyTMa/Kyh+zApgTl8DLZn85ks11jWxWx87NGt
M6xk7ig1QAdIa8T7SZtAiT+UoOC96gvYXQB6cb71RUkUHaumuQFT567npTizbQS6
mKLpl/1JCeUREtoBRuK6q22x62M4/TD3xtRTj7EWyfJuzMghPTPas8X1JpzBZ5fJ
CnliRsubi5xFTKfiaDiR/sR6ZOWkI/ZueTVlnUeHxsJkmQfLllKKWVRuLQp4PBLy
zdG+DnMIfKps9DX7V5RUA/gWAtBARR9c/AqWAi2OmretwYUveS9T6YLy5NKFQtph
BeKQMoydOWUEvnAYS5wwPgpzeNKj4qVaqXL50ZKxiQjme4jf7DyIqRdmsA/LFEV3
3fBRu/L7r/n7iq/irMKXMdgIp9TD9Bi9EzvLE9MmFuM7Ws92iZG7QY7i8OXJwBEy
+43H4xPfCzampXgOjXh6geNom1jOuwyLnP2B2wtlauFspEsZM5adr7sQn5O/vDd9
dcQUphzj195ATzf2XwoXJbhF9rdk+1mJZ/oyATHcTBoa07Euim6izIqL9PJLyk5T
SP8pDX0LaDIAmW2glkIuu5ciVmwtqKooK8merokTWf9upJ6Yd89xXzaWseap5ohC
KMqpfSAdCzdX1pEC1aEyDgrVUbJ518mQWgsrJdUiSgTxe8lnTvYmGjyCr5N9RIBG
C7XKR/SAVzQl9CKnsC+Ych4OqqAvJrAS40/pB0H6AzslascNAT/sSct7fICIXJna
sJoNIYGIId3HEd+fEF6XYO0P0qEJC2rquToT59yIl5TeCx7c4qI1WNjyHId5SM1J
lZedyGUESYQZTEImNCLCvoCnttUPvMWiA15ZTNcaJ/28aE+rFW9aZ3jajLbAz729
vLDNxBfjf04l5kwFfaqq84S0/9k/Ro2Jnbvas1Uf0ObguYQahQnt46JtxCA7+QGl
c7v5UkunE47IHZOO1pxPbkqD67LxDOId9vvA7y4dBaz+W5FQ5TYrfDNaV+wUvQfx
FAwnO/xmAhSWOTuak0CPOYyuGbyFzriiYoMkHdl3YakVdRpGcYkUyL7UHnt2DbgN
Gd8oNKH/E/5M8Fz/q79AH1IU/j3gGKd+IU+tRqGm+9Yy3UaTJCugyiTPVPXxTYuO
sjehhTIP4vVqqe/OqhJFlsNz1wU4h+cwoigXvmVAxNG7qQkHHoJ5Xy1t4JQ/lF0C
qXT8j4hyVw5hRGQquWWguTGkNVAsthS8Y4MBnEJZoF/3umX7a3fUHU/POiTLXO4p
Iqok7nkUQ83uLKsU3h4Ib9v4LOigMAyPq/gfoFeGFeJ3aqMhuUKumQZALyFhAs78
A8oo3czg1XmiJJOa9x1gv74o4bdXt/qHNHsC4mJ1kz/j6ZUjllkqNjl8uos3RzWx
MAhANH2TqE8CRYk0Snr3rIXlLNyaGp2jyVvk0topz1K0n0GDzv8leb73wdy3BG0Q
TANdEd+GCxS0fYoXSTxEEON8DmCHra/BUzHaS+dm3gpf9soNJI6AC4+nk0SKrmVY
k4ASRh8SQ9I7vJNm2Tj1mnx5T3DDIw+1ke3jSWn3Kd3coElCV+ORUwUcvgf8LSs5
3mtFVhEfapy0TgLjNGcZHyKYWb9pZdXG4aQASdbp60xCtOCbEkwN9hePtyXcWEAz
uBHqWtFz1zaKH8bLGoj5NgU+2suGcLheO6wjLjYIGKX+FAoSEL4WXZ66N+tqeTfo
Nn71isiVU8GwjwZCEhIgHiHPLYtawTxayq9oPshuHemAYvhHKPUS8euJJWIUjxx6
dKK7hEYNhVKgH0QVDLxgM8FRwhz4oFplk5No1VC3uI57QFdq9JPbRra3z+AbeUQX
lz6Kw/slj3LGlwoL/oP7+O1wJzarALJ337Jj5BeQhoPFMU7+Vj/SBFrVeOZgeTnd
ORIYGaTD95oEJhU6gq7EoieU0Xubw4/DOusRxkiQ6lcWbR/cCekTzjvby0bBMP0V
v2X7OrB8FgqUqIaExm/G7NQLtB9sttulFQgk0ix2d466l/Gb4VeqNpfc4DAySg30
8bFrQWfyNkCIGNwDw8LI1mDrWb9zEMpI6ncDoyZ7SaipVQK4b2nmGsolB0VNTg10
hv3TjN26ihJ4YwwmvWnOrUKC9medTq6qOleqKpWsNvkyXIJTMwViidtn2J79Ps1Z
gHcWbuMfRWicIdkA6VhbTvopaSZDF/DjLsrfAMSwc3cMFon8tJ/iq8UQZV+Xu+KV
FzOZaeFW7bV33O/YaPTXYBobScrd2gbjFyy67zLKKuDlCrlr10DWwf1xOEz650P/
2qROiHLfuzkWBz2h0gZTEkXhoph9i9nPmrIK73iyJKG4Mbm605rS7ftbyyzBwOPg
rd9a6ISvEm1PPYxU/oChgL8vSTGySRFg5JxVG3Fj8uieeS1JenMD6Rs5mBIoqZCU
IlnchudNz6HK91dZRoMGPJWt7lCN1V1BXnaZvd8wSeCNzukDkvAmP+xSNMM0ePo8
gIO9Zt/iT8GZzaUqnsnPL74ct4Ywc83XYwwRH2URiDTWHKVPnSCbRLjQfJdkEC5M
wvNJX/CVxPPybzjt008QSe+OFvew6vq6i4JS7sO7zok4N4XZ6gRvRmF30QBUwFvm
Irnt6wWuu8iTDWXF4lV7boqFFIlcMP2bgB2taYcBttYctmjCdTVPCvxp1EsKhUBn
w5pOB/IEWrONeUF+Xb7xPZ9Fz8SOM/59HH5q4ga0LI8jL6UtrAkZVqqSeCwfu5kg
F2IIgDiQnejmz+qDTVAD7BdCUo1BdZGEeK0QXEk4qMo7yZP44isGhrZeRjeyMgJ2
xKgSUj3RiYllmSfWCP8Ewm8U6pp3DrXnF87qxoz4RefSYxG0oyZgGMRaPxJfeZC3
F96Na3LJz1h7rruxVOq+AnmVGGXg1mS2+8wV05z9GFFWbTMBKx8xK2B2m/+oIalV
sxpiAwTBKCRaUCOiSDzdxpN2Ye9ff7l9H8J3PmLab9NNKPRkKDxi3oX3axBRPMxl
kUuGLlVR/AUKoyCCeBsU1FKIcGdJPFheXzpeWd5G+Z7os26FAiBNXKoYELTh3cV0
u3W8VNyZYMm84G2F0fCey0+l9gP+ZdVhEI9qgngKC9p+k3BzcDb6TLN0Dky7xqUy
89+VGiS1kgiQ/2X7eQAt57FzlqJI+Nj60FXqHixlO5b+CBDDaHg2vJDyn2ZuJaXu
kZdm8Vxx4JKhzvsz8Rac50ZJDB0TG3NlrUSV2c0P3yPR4KghZASF2E2Ax4rsghO4
uqMGMB5efZwIR3mE52iL1eY0l3E7LBZ/sViu/R6aeckJf3NSzan0NMwRtBes1NG6
ngwTX1VuvpheUAgo5OTJSK86dybBjRrucL32nKEPeMOyuxMNFddegA6IMuZPrngF
f5giTgeJxwk/9lUI2btauwCvu2lxVCwW9+VSCG7Le2dFWSsf04swo28kn+79PlkP
Ti22+yPMVm4ZBQtOmTRO0MMK31r5hFj3tFVGrWjsB3Pt0jLACkJ+/hu6NYedcjcr
3V4RqTD+6AWDQn/ReTN11OEKz29RUZJJlBrer4c6XBC5HQGdgmFvH8GQo81daLDO
5JqyVFM7wOjvUvxn1xKBQNU5sXIWvIfr0FJv4MY8cFvuvZ7CJxQipAZ5H0X8/y6D
7DN6b8eHoNUD+qWcI8EBMhAMNWEZpZrJXTAO4y8TV6Yv0A6G8VVs8TTFtxOAQ+jm
Jo1AfSzMv5RmkUKaUSbeXygZceMVXXYrIFw2CpCDuMAH3tZUBTN+8FLtlHQ+06SA
WyfjbxGnvyAc0jToLmLfKkQlCgCUmeRkTHg3OceILXtoUKHEcnIlMzz/XJVuWOYo
prfPnumuW0bHm+hU7JdEluabF3fFS/K6rQj+mDH8gSjwUzooeLfyVOdIOdjj9cmq
eFxgCs1KwDrO0qIwmIXclhpgR4H4uQ248qpFRWKRlYzZXATd95n+9Lv3YFDaNNr+
8a2+Z5z8Eu4VH0Kj3DtbkjfJPjvOPdBPcLDRAU9J9qYbw0rZgBirrS54kSX+pjW4
4lodfwgWGjLkG/ajdljw0Xl1xmhtb8cyjWkZWTOSWxW1hf6AN29GPlad1T/oYoig
k0lAObqoLjd/jslrnC+7o7s40YYVyv9OA/Bwo267MPBebRreHLCLUTtyc6foo66z
dLFQs8suOasZivKwcrn2qmi6Zz0D67FwSu7N66FzIbeURKhsNDWZ1S68FHDwtwQ+
XlqP5ZCol9zLNt3pjWPNSjP/wOv0lGpuyLsvDIwfZILv8YQ1RdARnQWBtTAMrUzD
cucW5BHNGnax7X8k6WVnPSaOIhWW6AkXBM1Kpv4nOjHonDWO47+TRZJC9r85iqDn
/pzRId9rCvd0B6VLpXpJI6hDdMZjNBJJE4baNh+cc6jE0TQxYzQPB5yhsTRG0+y6
94tVkcIM21K6IPREMklDXngZ9h/ikjpKgk21zVNUqudFYnXNTTaRkOUtpQUW3UMD
019bwp9J0K8LGB75e2tX8KaEw8EMCu5FRuSY1FOx7ockGWDaQKGJl+Hte3AovCXE
KzSNDWrW1/t+OW0L+KNm3NVSh1Yw/hpyi7sMTnN0owsiNRPmPocEq0CU1rE3gOMN
075n6YrhX15rS3TI6WJZgost49D8bjilyrtFsyw1M8nH2GJFo4q2u78v16rAAuCB
pKWgHbljV+M1CWnvEc/oR8+s0H1EF5hcdzVjXwpukSZJzXW3MAvB0xYoYwAjrhtz
p6K5Z8smh90LA0j9yaE/uBNt54knfKjKU+gFG9UnZN8q/7qQf2d1+eWzgMihohYj
StH9rdtlq7wPe8h6QR52NYe4JAHEcfCeMAGlVqclNPQjBq2BiTWFZHLEL/r3OgT9
TB3NwcjF2RvUCIEWaq2rrYY2hs2rom4Nn/1f4T+9s+qkRp8fl5JTawTglelbu37U
nEjZE+OY2O8dbnnGASi9UFCuaWp8XKwBacYd7oZ6PObhtFeQCq/AUSLpXKDYbFKC
aLbbHmH0p3pJctNu/XRpssptgv12tKT0AUAqvUCJSH4ty4pDX8uxKoIUUFVoXNcC
MddBYbhphpIy9VvBWizKE6j8JeIWOHoKMV2FM+YM1Uu1ZHV8YiRkD5R44zhEgBh6
J0RdNm3bTNgeeyH0KKGjLI1UlzrmOSPruAPvpC3+y+JlTdakmOCQFLJSJj3SzvCK
DXE6D9dwSkZTWneP/sBbLkDDZn+z6SwzbvsDQj0podvvzUjPCvm+T34VTp3n+uZH
N/qngNpIyRWFJykuy1BPGwxk+CSj1KKZ/SwsKr1sjS1BrVrB4hYU0r3NzD+MV6sM
UYXmyG7JX20gqWzBzH42cFwkBaDxKsg5zpY/nyYRLbEefnZqXkJxEU1lfU+5YFxD
wqiyRaCfKsbZ+pP2gfBF8NOCw2ZkeYTDtqlHpUNKAw8zkucCm8qZbSnNbm0PEwJ5
K+vWc4v8j+pSGuSHtC9TvyEf/evCN1wbmeC8gdOLUl4le3zd9/i2Of8lS64pIIRK
BRfrH8xvXjZfqzMdWXvpUN+/NooDkcWmtwKSjk0sQx3/7InLEH0DEHTEnYBv+ew8
DEp0+5GeBRtH0Ad59mLX0iEOC6THPc/NirHZxOFRuePExrEe8NrpDoPs5I3wLaz2
Iwxf+GkF3oK1i4eW8Mv+EnqRBjHV2NGNxtkX1r0mO9EoWsijgYEa9Ttm1XFhmmrv
c5K0vob9Q1eJgeZwsy2moi4kkNGoAItN582lnPCZV1DfXB0v4dKN1h6wihN6dJ+F
w0W7DRphhw4p2EBI/5eGOeqQKXcPDXR0r67jE2URgv+HzoTwDW1nkUH93LRqHKdX
LCPcUtWChYznETcu7/+Z2lVzohzjMtREXBDgoNMAc1ey/1YkJrujbLedFty37+Tx
LS5NNI4tdvH2g6Dw2hEKk1MCoDfe4vU0+WgEJ9YmqMO6zyp6/tpsF297HTeFd7qk
XIX9IQfWBaOauo6TgKj98ToE2Xdh/xInSDval0WQdQJvCamShgPs3A8u2za3PBL8
E+ieCyxcF1tosjW3GrVh77EYJLXvXD2D4a/U2H8B4zMeMnN22xW0ADprfYbX5Nb9
hAjidZmBAxSnWepZRS/IblBC4IAY+O6zc66p5NzxBL7AIZoL3REAnep4LHj2Ce0t
hj9RTZiWbV+LDrVZoCTJ93X6Pm+Kn480HOh9ygd4NSOo2ZkGgyR00F8tp2guxngd
83tdzotGx+pekaPtbadSLYgej5DMGBiPmc5uIpm97f9kteq07k0M1i86d5Oyh58y
3koksQzGu5Ub7WyB7Z0ioBxHHNnM2UwaMLiZNCUV5hYbeHLHioiv07hfwqFhxbcf
EVUSJgd2XKkViVdpIjlPkLiFe9BsQfQn15cImt16wVT1+C6CDqf1TgUdltyH++ZU
ZRluCuZT8KPOI7kosVLXVMQ1+gr1D0EkFt4/JgvPLnmGIc1cWpQaOKetdZ4KDwR1
vJFoYyqShWTewZwWxqqyaSD8D37yEpxPw806/Yoe2NtTyOq8jZBDAp9RkfN2Fp7/
q5IRa2ZrC3JBE4CvTHqxt6oBZPScj9VGsS/cCPu3Ljaj+N3rWvjFIK3KHSmc8ao8
2+LQlT860mV1x614TepGovCURRwcWHv9stnUJQT8j8BUsnno/AYFRM06s9Alew9i
A38jstbcrASt79EhFYNf+X3npqWeH+ScqcsfjzqXyh0xIUnAYcVrSSXQo7sVg/Ij
tCOK32rvTf402c3P38dLr2GbHo+tewUc/E62R3mxjUmgfwBeuUw8JNAfzwCJ8wqt
HforGKxJNMNS6x7ixoFzyZRh75NBlUnbEZjJ8T3PiMdrl5rl1Y8Sv4N9SejpdDnl
DhzbFFFTn8nYqoibmUpiwsocOyJawskEnaLwjEA6D6osPO1Otx8FMfhukxv20gCu
IQTeCC8BbAprG9HwQQsJHO9FgnuI/P991i2E5exW/nkbeKP5iRjfKtkhHnN2dgbU
GxbAq1yfpavd1SqyLZLCMlVBHNMz0fO4I2GcuP70Aw7OYFQE7rnANKqzfJ4f9Amu
80qck9/3XL9WxiM9uS8FAeP6msxEZqBmBmyn1lpF6w7JM5dRfWuN+M39AxIr5I7M
dWh7FfQWTl4PHdHCanUW3+6P2i0CzFUBIA7KKakvqEbITLGMCkl2Uh6wXeOmpFrz
jw9Ac/90NmYKWeg+MLLW7R1+msIeDjGdB9D8bg4cNlCzAgyCh6xmCQgCEoWexGlM
dfNTg/rObAzQ69Db2zWtG6FrM9ZlK1EHcSH5PqbdtAIkpqklBP+ICN8Oq2a2fmJo
TOtnuAsJUyexGyf7QVyxJyuRbeoVG0dBVSLS7eF5IdQGEXaXxHI302zXOzp7h50U
leSiHi9uv86YZ0CYUMk3U0oUMOOhAcH2n5fBr4iKMDoDZGdBYoEzSpiA7K4SqJqf
PitZMYF13kClR9hwxvMWAvOToATcDrcRqSUjT3Vu0AH0HdHcSdCvesG4oNJ2KGzL
hxUtK/ob07DaftWgHAdd/eZvTD29O9UczTDTyN7Z6+WIP5mTxaka4VqSm0//etDm
rK9+c2NCXgZRfE7xhjREZLFhglSaiYW5AGxnnyM1IEagAgbrat2NSWceVd8McEjr
3WwQsFofp8thZ4+LV5EPvwgw9NTsRwjAaT50ZaRugpvpTlZgkoCJYpBXUEMpdmcP
wsO3nBuFwZ2kaXhZ+XWuPVoYpUQtFrrqqnA23Nlee8Qaw1HdexJzuMUxDzKOUGpg
iVA/p4eBMnxoicW7+lRpYL+VTr2NgKQyTCTdacuETG/JQ4WaUThfMV2wmdcByxjv
pD9soe03mvVbCHyP5boDiJWqkUShW5ZyVFL/xqyAgankOPO+e/ZcdeMlQ635qun9
q6LgwtfX3rFgSpBOjj+NvsU3HXPNY5RIVo/DD4BKGT0q0J1F8qFIrE4t+LVFo8mS
aj6/upNKMFw7nyd8cwpe+rtKQstP49JQiL7KKAkQPm2JulbSO9TAY9A1oZzpRU8l
RvqMQfn9uILlI1XaWHnhJCKojxM3FmdmTDnPvsgyPQSoCQZBUZmnNGIQALt1J6ZS
MomruN5lgkfOC9FKRTQzuA9QRjC2te6V0noKufDnuZecFv6RTzK70iUjky9aTOef
iZQf4X5cLiIdMPwz3emy0715LlQYwCTyay9tJ1oCK/KMvwLD2KSLIM5smukCMFuU
TguzyQJb71Jfjxel0n3GNnYOwJibyZD2UurTyo/a8NYMC4SAIETiVMg1dxJm2TSM
hYWgWJj97AF8zizzfuzTkNmLKfEC1qAuWWBiQaSp1rpi5tWQYqdC0onoWNi6lVt2
4Bp0OLRenE/7L3Nwq3qr3oBIIk1V7dpl7WrIzAwRZR2vVM8J99+Ox8vZaVDSwJg+
gog7aaOIaUJhp4hZxEm3+bwdGkGjZc1Wum9sfOXtzyn+Dc9vQltM1VI1Ute1gK65
pb19mbUvXX5rEb37/zcOogTlKpZ8KGqvRYNQ2f8m9zO2CZrnmkmK1Oo7Ytv8uJ/k
X6i0Dxem5O2DSaZffMemeEH6jMyAXmLbFVPwJqEtIcmdGDA+YBF+TVf6y+Y1+FXV
21m2rD1q8S+fxElYP8qt8dW5Dk9Xp6+HRdQ85nOO1ALz90jCYB2NMVvvn1s2g+hh
WCdu8HT+h4d/cconLfZc6THcMhzBl/wQtkA3TXSGYoCyxkMf8E0xJo8hQV6Ajrjz
93vPHm8dccJcLyJBpWTqZy5jV10ZRcB6QPznVICwmRl+wvBY3IqCoprpWtuRD1Bl
A4jUj70+VFvdAjUWfT8MFYtKx7myTkgRPcXFQRzduwbJ5wEyWD4ANjS981jK74sY
H+UXDqmIGanNMOvu1vJKUCAyChOk4NH/Nc41G0X1ITkbZh1hAvN65KKLrTQ5WI0K
w6fz1BFwjFHgO+gnypanHTmB+ZbnOk+DljWgLJhuHHrC/3NBHatX1k8INcp6htEW
cus6RmVCMaq7cPjGlxzd/RguUyonRSADM/KinIDdflcEn2egdw2offgBGJOGGqZD
+8r85CMFcyEUauVhPSRzX/pa5+Zsmd1/KNqesxrLzGcC9nCU8KfqQBY6y4+F3Kgm
QF0H+zsIr2yhCjLNBJBT0Yd5ZKNpk6ZB/gRImt9hGQp3Pjj6KkxNbfaalrw3um6q
Yt/knmhuOF8iYmd5DykUMWkQHfpZDOoWhXMMV5VXllXa6FcvAKjbs0JQ12og8obg
Zl84KMPeu8nSCKnFFZwKebvZxon6qqOTTf3PxibBWGv9L6KsHi3j5OMkex+Q2/v0
vaid9v43ZBympEId7s7TzPdS7sWNbZ4Ds5aAUPNyFERA/Yms07lVJlD+9POKKAS4
ea1WSWirOErfRSv7CpHkyDTABhxDPZ054il4czx7ZqwV8luULIwBqkRhIEAnYw9c
tecSJY0lKtIEQaQBw4Y2ZlPr29FLzRwC5hkFqKwdMt9NW6voJEz+f9dSnQEQUHfN
R8a2jOgiFJj2UVEb6e4rYIytBy9UMHb/bblDBVi8199tsILFOtOGGMWnaxbVx2Xc
v9CJwJIVOq2k10IH27i69+Fc96u9m2t6K/D+LhjPwLquLr4j0wSJnfJw/HYBxIqT
LrzflOVJQhuGCVXPxiCoAsZRY1IMt3UaMt4QAPtX43R+h9mbapeQ2MC1q4iRXK0t
zAW8tBlIndaU/M1QOmlOhvkxesauMkz/Q9ZROjhDRlO0sMJdIJsUJHIVIA/K6/7v
F2DPKXTmQNUn2zjqfN4KUtxzVPIJ/NnJ0Cz2AipISpMgVzlxQMM1CU9vqfmnVA2l
UfsT3DYb/5QGRR+W75616TcxE3DUgAVeSsIOd+kb9+LBhIEDpLUAK1sLwqQa22SI
KOJQ/7RXT0vJ27/xicGCmAoEjrbyatqfgSAoE5oOKSOKDc1ulJewsAOz8DMcF2ki
LdERMNynpL+lm81jo7TbxVvaVB9ib/YEtUUmjDFMezkbYlfbZD9GqR56Gs7CU9uU
e/i7HO7q5MJwo2iujAezIAnVQwnKp+oNhHOp78CVw3kbqAdzItHsNZNjkNPM+atR
KXefb433I3gohKPbSLYaal+owl8un08fkLTs+J/8l1qxMLu+C0IlhC+cKAzPjU1z
PoJ9n/WfvCJPBLt0P7VZwaVt3e2GAwTw8CZqbNNS2iFYlowCsoUCrE8e/ZUDlAec
3KBCOg1X/Ur+FxZDAUxtITPGbYSnklElg9SMewZGF1BJ0DniFzOpXrmVCNhTj9O8
jFlxbBoLNIKh2PtU9Nfkb2wYc7zrPrHkvFPjKv6rckQYw+kzPqbDB9Njf8tEm9T1
1V9B5MQ1dnvGbqb7FJJDqZFQBs3JnvPnfyVgS1LoMwQNGdzQP1LbQa+uJ5qnuYeM
8pG3gvi9Zqhw5EeyPgbDcxIH7+3DzjoQU9AJ5ozImWThIP7iJumVwss2Aobs4q+c
UXwPC0SrUJZgKyfckqRBs8MaT3v7ku4flELPOOgnxtRqdP283DI/YMn+msR6/NyX
s8bMF/6DlqCQqRDFjLYpXBYZQialAyAKDr83xQlZz5jfBusYP8poRdo0qpiGSLyt
hCFzPAMs0r++qM3N8DWVteAVheriuI2ps52FfmL6yFEjpwqY5D2A4xnuL2qG7XrJ
xvwOK6rVlInXMkJNyi2H77w2QRWI89wbnhv1hs7VOGw3T9KUF+KR+2ri/YLcrHqw
mjzcNL72hlEyVG8dlRfCgT081dmsE2AhsK3hgPxx/coSDtt3FRtlvuyVUlV464dL
sb6YaeOGhTNsQwnbhXR9CaI4lcsOIUhCdvplj7WTkE73xmT8qY4HyITiAJ6tR7lJ
pP6Gu7lUgEa+frpIQqI0Ty+w3+73DZ+yEDmA9bSmqwFeiV6oYQYaXXFkgnV12GaK
oHXinBMipSum2ujBdCy60HWo4RR+EaUh4ocphXXyxvscraz1EvFgrmLdG8Pde8+x
x0we6O2zFF3Ao5TED22fGA359E+oYwc0MJPS4+C/L+RfejTldkCbO30asSwOU9K6
DXSivQK52cJWu5X7AVjgbqANj39QM5JpdxGpwuPjN9ccVKQDq46YsMuLSMP9S/xs
PjyXdxqyO4D21vSRRah4lnYfYf5kdHrdD5etyEEj1eZYeZiJm/69xlwyvZ7gwERN
t0+fQ1MXSVyhzDC8Rfe4etMwBEoIWkTaXUS5jtJOk2TqtW/Yu/E85URXTCSGToGj
P8W/4F9RhuPZbtsn/gQMdnwy8z3Oo+hADsJpN+03j/MfNcPwU1T32Axm3XLUa32e
8iRBpbbZV1C1L/ZI+QmjV+hkYTUIDool0hw6R+jbrRIbEke/SecrZwiTkBs4fzdU
6Fk+Nwi6J1lIZr/ZvXiQcqx9JqrHxHUEGfFybfWhuAfviQ+upIGdxEghbChUr+Wg
CYnt8fEH7SaBDCO/gFoSHnBgqpZXG0bp5EsJeeZpJC8lKFPl/fhlsUuu5JX+WRUe
0SQFsiMlbKK7HNVlCX+RsouTIBog6pDSN61QQRS5g2OMVhNo/MyyTOVOWNlpsGVi
7oqobAT9G7dVTOMScfzEZTilA9ks6nEBuKdUIc+oNVKVQl197Pe4kRAjghKFaRee
jNGLRNr5hYj7olX+Y/EB2eehAxsdbs3LZODKyZIdXRsf+Bn74VkjDfIMR6T7dTiH
tlmP56DLHHEfcGac6vMWfuGoHrD7OgzcsnE9N3i+T8dr3s/UCPqizjekN3rf0koF
gl+/0KN3q4rc1lGf/EGWk7PhKzIgKD1IcNJGb0OdX70887uVLa7lrUz9+moSnWTk
tF2poXmqJhBFlR5yccgCkxB+zTm9rocwUkGhlGCeikfbOb1FlrwdMsqAeEb+pfSM
7HptG553F2DXAtiHk7nfGtmr8NKaxNFzGv4jhdK5wE7GTZ1ZSvEX6GchaxjFtVXH
HXfvMkPTvwh16wDsW2QP4j3IOoQtn7OKzGhh12KJ0xEmOfGyyFs+5thC+0Z8fFsI
87cJHSCQTeb78VRCBK3dX2JIgoB2vP5AYHc1qAIBhJxQQIDDkhZZpZX61zA64nMT
sn16SKOptcYQ6zji+QND7VPFd00VgLoGvPaxg/1usRmASiJihRg24YL4uGIWLdDu
co25nAxkTwtJTJinlnLTqtVVDRlFDnmw3emS7PUQHvdGdzQvGNw/Q4csI8EQlbdE
h+7gDCQ5BpOPtoGt/u7C1oL4uDulz4nSafhbsNqVxzTIufWajWZKeW3caet7Fn9F
evaxyeso0jkZUlU2VjABo7cAIfpNRrSUikU5ZmCCi4ctZHSN8UMWMsikES9c33ht
2WmVhz3JyeGvMx8HS1SNYGZNWH6KOwwpcffb8kgiAhUMZVx2cn3m3GUBBgL9x0Ax
kM+gChaHAnuiH3piWCtKFJbQyGIvceNNDY21Fl79oWpmzP3LXb4v8y8AY6IqCRk6
t+Hf7gj4cVT9aJK55q6ZD3RwUz3yIx9wAOCMp6kf1Di8oL7O8qvhGKBwn1kEsE3h
E/iz3jSVjmjOx4F4kc+2Hz2XS+AeMizF4vONhmNXNKIDqKAVNpel9e9XK93pTj8o
grT9lKV48uPDM8TUKxW1VJMM1LjPbK/OqQ99ktDyrn/HJsIiMgnuV1eAv2thW1we
ukJ2QYB75Oet1Wc5QfYzyFRjKiJMe6EcFDwD6WRMO+ChVVR4RAreJPHrAt08gr3d
a5BcQuGnWQuU92bcCnwo+iUBVeoh7wFQTZo36D3lRjLw9R0ra8rSdtH8NbhkiSF5
ls6BB/mc5/KWbSJMsL3oYkBltTRGjY7VMS+B9aAAN9pMF1iJyxBJXjmToXsqoAVV
Yu6EvjPA2fFYCBs7bsk6YC9kG0mYotzYXWM7uUYSnsn8l97vMoLF1EaK7hHPvoRy
KN0qGBCOnvJRqVRjZSO9szjzSrdg2/8T7qWDrgGrZjLH01Afe1vtz6UzdKkxk1PS
/vm8hseqTd7zdAKhzqKjwKVfqNOvcGiweL/BPlj3Ju0eHBp7U72uYma1MYS4fkfq
te/G3PktX6cWdQvH4jdjja+Wyh96rdzmlxfJEq3V3BNrAEs6aZzP1rbnnbjyFPQ5
g9bqkP1wLaCrnB+MhbwRriyX64fi+vHWkTUONtfrQ6B4/Hj71tLdFZNoCus4Mfwf
aWsgJ3MKZy5UWzr9LDC7AmVLNYsjLO9LxGg0yYpINpvrJoMDsY3v5otCjMAkZPFD
ELyiyT/cnqWAHvsTu78WKhjB0J8MTMp2BspITD6p3DUjpC0Cn5eIY+YPZqLtXgOC
JQsIssD8S+wcyHKPYnG5jCYCz9Aht2X/bGnmbVGNCUEdy3XLsP0vmc8ZzeYLHJwB
0APSjbP53NQ7QXuYf6T0yGil8HbkGxMnVoyNMfi6jjYHZsLkz/zLc1aiyFr4qC8W
Pp6mRUg7YhEnch4ofz1XSzSpETn0yl0lXjxcfZSNQrBEiflR7b6+QrlUViM9Qz/J
snTvwk5Gy0KNOcgekYLSgBqWL7WG3N75o6hBAoMPAw48yFr9E4nqZZOBpu5ioaqe
XG2KBF7zCIALpQEDVA4AyhfgcjfhZiR8xPn3p0YqQh1uF0roVRvyqyCCJ1rIfHAW
xO89IbuN5+MVZLUzJnKkPdYKE615KtFBGcfIXKuR+ew4ww68gxsGZjF+BYaWIjAX
D9VPaPHl6+VV/LXDwX7/brmdpX7lrXvCinxRXjBpfq84PWeRYCSjG2b7dTcmRQ8p
3bS5pMlyC1o6jXKPwl7WlnRoz1JdIB88AeNT82s97/EzcslFnmpPH8/3io1l6K1S
zPsJ+Gd4WG4ImZUI+boZXOj23BHrQo0HlLqKSOTDzxOV2KKvf0p9rcyzssotjqay
WPubo0CHwCWFp64XoL6m80xPCwGrDPs2m7HtAVsipzQSNU3tr7xN+jx2AK9e/aH4
bQ+t6f5CGqTbK8Y4SWq11Cl8EmKQRY1i8kJ0lK0274H9MPkBRKibmVKouFJ7ml5R
5mNcN3id68k54/eJNVIaNS7sAruCl2LGHlt3r0sr1yCnD/b4yuBlQ9/a90Mjcp4S
5+Ek6520ZAdJkuExz0D5zkBLHs8uE4FfM22YOICLa7LxRUxt+5/j2NIm222KXKEk
0GJX+y3NdI2UWLuEgsufIt3DJ7uPxsT9VGO/8Xvgw8/zx6Zy4h8DUNEylTjRecw5
fPn0iugQt6ok/W/HLkafFjcMMGZpekO/vvRPEZoBRZEOL/8u+Fk7uSGMYScdJ1WV
l09fJmLhqOjj9xQN/A1ymgrD295afgesnj1AV4+fovpPUiqGhrPzUVTysBUFkCd+
tnR7e5NHaC4NiBbdV0RpSa8fQ8pVA4WRVSCaQy/3dPKrvYjBG+ImJPhDcODtQfLn
f9bcPnsjBzHzhCGw1/r4v99J8hrjT8tfnkJs6B+MWmDCojSrIYzTIM/Uk+24jGcn
zqyDlWgQMGx7I8E0Rs9zDD887rdDs2ymtVQqwChCPDXgQ5LmTnN8sa6UcSwPk7an
A4BjK9WGCNC+rETETJ3pxLQ15iK7kbhZoa+0e7dzt9WjHEXQTsw8yHFw89IgH21i
VxcjE4c6n+rVqsKUmU1mTZTjfo9qbofB3b42Q8k7dDNeewm6x7UhurtfjTpWfylK
AnTUKvYtOY5IMivIXaTszLw/LCkjt4r2aznVzh+iE4iTPCyijj/yhU8JDdNg9NFe
2e/HLK0DR7aJHz8Tk3PznZF5WgfcXaVV2MkpUWBE/z26L0pEcDpea+bHzF8v21QX
8djhY7hSbAh+qR1XNV8IWoPFanaNF2r5qeK9fHGHd5VmRiny6tkEzAjakyBu30JD
MQT7ig40Jqfpd5dJC5GkHxU8GBJrqAzSi+QshKXlDxDS5RkZnshdrsJPB+cS7Bu8
0tEzqKqnWgi793YzapWYvJSo8ESDsl/16wZYw+tB4Do+33sq6sG8LnFJkt6kH9+Z
Qwiwx4JJ3uqsx1Y9hVih3rWVLMgEt7KRJRPzHgxqOS3Og6IxFUXrqAtnoy6GI7Rz
JgzBoWgO8Hfmc5X2dkIgK9ljKVgc1qTjKIze/12EPMz3SQfj3BiaV0659WGk/teO
ZqL1rTkE33LszgsQQ67KjpGWGFYpgjan9BlI76xz2mUBJ4nIpTUAs/zpgvE8Jz5U
N9y/O9nNyRxXkdxTcGJWg7m9HADhUkn8sV1pALX7Kf9uDoKqNHpKbfLK5LMcJcY7
0K86Y86xXcjaUtoV4MrIWs2PUTlZGK4/7PqRIpsFcro2tcsdkcjvuWv36l2xq+ut
oHk0904tl54raghTa3Fbv23Rw9YF4Vvbetz7NgzTrnSBoiDD3n5/Q5elSNqKDCgn
9CVk9fLO4qJS+McardMCX/SOjYHTRRdQvc2iq2J1CxXHGJEFmKBBgcN5DmyjTGRq
+/ijn4xmTouZlULLKQbv8EAQegjsfl7s3Cs00Z93VFAlbvY0NzQjgoKHGEP4u5l4
1UANhEsov4bsyfq/WVBf07+u/AJw+fDbFur4ZE4H5dRqSaRTJjgkiphHFDIVYbcn
LVrgSmTlTHdw2aRmbG6axBbILh0aHdo1rDQurlcE75552IVfUQK1T7L+yn7EzJmn
XoEhMkhSCBzCFkPxBYiW1TQL0SNnTJ5djktlXOMVckxIKN90fn5H6vpyNk+EBCNJ
X5278Fx2WQOjmTy9sKU/4OC9NibGaZ0EQx5CmunMB02yVgS8OXrqx75mUn4omDjz
mPxoyCvliVfLFUqjok40JOx+CLILvK/UbuVzxv8iXoH9vUZEaQ2z5FUQD1qaJW+P
tdA/0hNbNN0CTDop7h4PeQDZRX+Fv1GaeR+Lo1QuPQ6cffHjZAHih0iLTkZoEHwy
ZRb2U9guonWyUHN5AEfwoaRzdyMuStSqCYens88Ap8YmToB9iiRIIw2I+ZJgppM7
JCcGZKmAKdeiES4QJ+Am16Kd19t3WBZCJIgdT5veNzIIhneL/hh9BVsc3TnYLEDE
M7OmV6V6BLWqxw2HYX47YxquvrBqfUaQXtw1AquyKXRwCe8CyyKMu2L6N6/rGUd0
xtp7oCs2fTZ7Qdeedcbh28BGCZqDJLA8CBIUwheXwzjUbW4vN8ounuI1+jNA6h+j
0NOJthFsb04T+g6PeWndqVNTbM1rMKPfXTcw/jMVpmFQLsHv2Hk3zJJCGzkbZKBl
7nseCnxkfh2ybSmjFQcKeaxtRwy31n8qf5ZDfqGTzQcDWBNShoQ3QCZm9ixtmHuc
kAa/cGEwx+mIbcS2BP7a8L8YS8Ob1cR0YSb3IJHsELLqgX1vLcRGCtkMpVvQk55F
Xm/SLV5KksvNI6T0r6P09odzaLdjZWQhMA4XEW20Lp4EMapvRZrpVR2miEcBg+yA
SLztuqAARzb2Yb+RKeaSUOjkUosIJEvaMcCVJuJM9KcBe3Nvj9dJ9m68kIj9Eclp
ezneAwvlH8bWf88qEcfY4cfgpZCZoREMJBySDyZQ1aWsjAuVDjJC3ykGHc9Ngmi7
3NMj3IG0VE++oNIqBCPSZZIUnDEP8ExcdVW3cuxF6i/f1kBySqMtEHf/CBMub+sJ
BMs5GPL4MCmFJDDCWPCCtz+CNtUM4p45+yK8GKs+vMK2ujFd0PFF9M2avsLD+Gdh
yx8QHWm78jFbtVT2efE6GIQbyAVbZdPOZmQ+EOzJWwy+rJxOriqNTtP3V/jLV9oO
NJiuVENuJwdDy8BVWNxWtNvGydIvmgXWoJtfMAKbUfhZJGLOBUS7nxjdEfIywru+
8LRwixPyx6J7w8A4zfnklMG/RqpPrKB2Ta2U7JrQDP6owrNO1l1WoBmzaQW89+aX
ShJG3BR3fkBvFdsDDP8hKQLnBUcOfv5RoKkqpuO5VR1AB593MQtjz6TC46hRWdZ8
2inA8EX2cYkZO+/rnAC1ULkQOULDFdpJJNXahqfYZcYU2u29ecWl1hKn0QCsVrZ6
X1ux2VpvBjH5as2Tck7PpB9Huxj1zmdR+tUy5/vHAHYAhXY0IPXe/SZro35pVSmK
RJDmy2FwkgODWGgCnoawWE4SCg1AtgGaLTMMZ/GcE37qLj/w7oQAOHXcKgowP8xd
nu08BTs+rU/m+Mez+mNjI/PHROhh/5PPcmRplmbpaeICXYIfQv0lqBkNGMQ3VJt8
KXQOI3MCjLqZjn3y8FS2pIXEkTyptLCmPBpBXJ8deJlMKpR3psSUf4Jf3SMX6YQZ
QWB6KuMD77imVCKeKZ8cn8VnHyqrXSIRJE5hNf/VfJPMH7RLNZEEe25olMjJnwzv
dl4RKTeWmBitaT9gK2Sdq4q5cmqgJF0JFBf4Qf28SJuNEGYIqhGAvnzwhIMlmP4R
lqMXJkRywoACLRxihgm1iO9blXxJr6KQfX0Q34zBWnIxwAKXE+DzSRwyqTZYljuU
Bi/O3jqlY14pRTQQVSfWfMjGdoP5dQ9fadbUbZyzsQA3I9cap5bi1Vs9I76Q+SJn
XrxughZHpnTXtwWDTI4ZCU/Yo01LPm8RghkWyx+6gVLUZ7gIdkkW9yC7D2burwwk
JOexVCw+xNAz80vGa4kaCZtxZOFZ4U6uBbE+xdc1X4H+qravOEP8NDSjOwLgQIvt
dVMrQbFmsIcBvYjM0x3fWUfHkJjClgS6rzJbS9ISVvFSQp98dWmUkF9dXPYdpEbr
Xj84sxVipmEBC4xF5jVwjR3c4/h9cO7C5UQmUjJ3ppzaizcPmQGxtg1KDRps/1h8
ToQO0bVhuEUtY/uVyInQ3hdA0nOHGNTH31XhN930w5xbYDihNB5qlva2a3H2SdQQ
c+bUb6Rpl+IcX1vkfNmqEMuncKkBBx9AaJKvwcqLpSLWDY751FNIrgF969AwB853
4PWv14MA7Ao2jefw+MEbPr9yG6p81UIl10r/DxuAcd6t8DNd6uqXyBI0XkU8jNGG
SaTrwS0q3RwUX8ZlIxK8n9P9OqBHIZ/MpcDiUy1Fxe3vPzSmEp2EiEfUaniNqaED
87SebRnz73EJhhUDOQ36WXZZFjrxBhs3y0dlgc3va0woxa4visz/OqR9tCGEEq5+
d/nm76V9rqDOHAVNwgTP5uZq3baU/n9uVeR4oXSOA/eRreSJhrff/tYfgjA1jVMV
w4qIMXxqnvI++6WvmvIkuQqDev98K71AudLLdFJ2fPlQKNdy/V2ywq01DQYiGD0g
+ylZEufKo7qGlDs6kHlthrXW9l81yaVYYVW/ySYqysPZMrLdBetifr4+XrRsK5mS
B86ziSjfoIPHM+sIDqXYIrW6KeChrMBigm19fXHZgTUGF0j2trGs3w6KcZxK6KuI
zZJu1pkZPlJA9z309457S9Fn0P7FkBP8srXrNHUwsFDoFkApHhoTEArsaaQtUE0H
jG2hJGTf2gYqFtN/BNZgqNllCzQB4HS1v3RUBTK8hqDvMu9hAo2+yTC/mnVd08hK
apQXY70iInUF/QfUPwyviWf1xBOc8mai+Q5JFVc+UBGJaoezB3aO5re+vJ3eBJ7o
/F5eLE8fDAILk2GiFAdk38gD4aoRVmKx49HA+ST1yKZN1mNz+oZyLrgVvHpm1MJd
klbf5B35F7HOxz8W5Ndq7gslDyESboW1XcfXikpnTiTuwDWFWVaiT2n2OToH9zZ1
zeeiWwSHW2X/gEa9y1ClsvrzQydkD8cug0lavU5mMHhi/PLNnUtsrb8eojh55c5+
DfZ8muS8Ro7fSY3OeI65IPEnO9a+Nw6KmR5bd4cPX7Jmw336IojOm7JIYOUqy3bA
yYkR7emyJO0Ya+k29IO0m2GPQvyhQ4YMYh4AdWY4U8njIWpmRNzd22+MZuP0SrE/
kPPp/5PuwFegEHHL+fvoxXMmWCRh84BMSPgmoLJN1TgEVL2n3kqTeVrqp1rTQLSG
V21H172q4jQIlx2ra8TCsoD1Bt38t88ok9RoSweTAg1i7o/RTPunJ644jDlWWsas
1Pq2jIFq/lCGBwxlvml97ZVBc9C+ltn/nvupNz8fkE5gQqnbyIwwoNztDHlOlCgh
XuANGX6pB+7Z/5msJrzAx8y1EgwC6Tld5Vx/xQ357etUy7VZsWj9EnPoBnPhv0Iw
wl9LWS8ipjUtOv3/x1MLH6+qYbjES5llkwkbIi/YjZnSwNy7eC8lREn64B7KlFS8
siUufiqhR5lhIF+hVFxlx9ERJ77plu56TA5AyvqVeHQeb2ZU+4giody6uhHGyrOs
+nuwNCdX53rpk7H/2KT6uEn1adzvBWQjRva0Ut0eMRsaitBzKYrZycAk+6smZkRg
a4pyuCL4AV+qjkf93W0dHsKHdN9UnmuRfFU+NHG8ShODuCEY5f8DQzeV/jTsr6KY
4gBjPUemzUQcR/ja7DrrnCWqxEzfy07IiG4kRReh5MX+3vHXoSBi2Hh6UCe3bj+D
qhAjYs3sPF5CF8Q1K+LnVZd/+dEAQjKJIC3Nzsdv5/OwpOnL529xQD6xF9lBGg1p
Nq7fiAmmWG7ujL39gJRQp21/4lDIOMOGKaeypEMEZXYo3Krznb0HOyLtsAKAd74J
F7eInDg7qvshehbN06YClFNuohtkr7dcfPqwGtSjsmJyHbRFZz/7TLApKiTG0bY1
tnYA6qUBLtH3svLWVe6WkGON1Q8aw8puAArpvYVAIiPck/GkjO68yT2G5TISBQGq
1lhoJ474G+mzMoEbINr7a8oGRzmIOJfWPKcKgJdJ78cu0cUCYpVLpXn5y8YaZ7YL
AtWPD0qDF/fPLlg4bg6TYxF8qj7V6NXFT+6ag78176lTCqzrLz5Rl/y47ljeceGg
GGmsOtz3ScMVuab0efzqhuf0K/YdDC8CMTBc9ZpV76racym+Qv8mu4IVlanlz89e
8PBIlNmOkLlMgwWcvj3CsPc+pIrNuKhL3qCXp1Frv8yqh24p7wpsJG1eUJch4AlD
ldS/KpwQb58ML9+eoV/Clv3YcKcEiic7+7VM4rYXey0+VQPpRu2gcfKlkPxseTFQ
9rMJVDrzE3Q4fu/6llmneMc2DxEoqhUob0gvOlgm9AhsudADMGjY/z30XpQtvbW7
jhKF8TkOdDNONxNLE+/zFwm6X/dTxAGxXS+JdyDIPxEvMn2PfuionxMKQ09qsmnR
u9/Kp3GgnujKeb3/gBr+nPtqQczzfyArWySAZQiGHJRAj9PGa9Pr+WFuhE9znnTT
PhatD7I2j/WUAuL99RKSEvMNsbigvejkLs5ii7JGUji9y6K/ST2RgW147Y4pw6Xu
iLZLIMU1V46GMaJEPHjikK3W+Zi1cF1cJPfA2fMyGyjCmMMGvaJcaykgokmF3+k0
wd7PFAAGEcvMSe2p/jZRmnY+kyCtJ7W5V+HinanRW+q6QOG3irCjaAyqC94l20Xw
Y5kdArBCX9VEEeN1noF6qvXB8JbBphBe3gg4NbmEDOmxczkhFCJ9bn2uzP4I656O
+lvC0m89uSNAIjHaWl9ExUBI6YxcjFIhia0KdowwsY/PxMjy/qb0macvKSXeoM57
tTWC9WPQnVR6wNdLVgjm7Oee0LpIKfMkD7Se0/K7hZc5Fcr/NePmV1X/7UaptL4u
rH4Zbq9aUPPSv6xY35PybRxhmCzWs0WtB36+V5m3Dup/y+gc0Uz6kVOhA64hvlfV
s7RlopU/QNJHEaLUjhyggrStgcaOxdjPXQ2qsELb078A+r692OrrA4apTU70l1y5
G2gHxgX3Pvql821Ffa0LCx3nuv08v/Waw/iWMzd3AZKN+JxsT+WJd4FNtKxlXjD0
sLNlC6rcA248G20/AodkSoQEDO2x11GxR5tmOBg6905A9+1067zIAPiSVjdR5SK0
GmombtyUgUakXIaEd4+5plz7do/OJcfjSqvXJOno/pIkgZ8Z5xaGqK4XywTNvVqQ
ePJcEt6MjohCvTwecpyiBvyQX3VhhW6J55ofur8qKv/IqRtlmcbA7mT0fFkFFQ1Q
0FGvrT7nRvb9VP0kHEF+Mkxw5ntCwhcWcB2XWj9IJLE7jfc+qpjymqWN2x4mwSl4
eK82J2KIDmGq4W/t+xXZJj1nSfgKXTVMs9uByT7sdJ13GWFL2ShfhS18VFXufMBA
MUNg+X1Fk5OviUeDc5u3hdaDGaLSzOt9jGTzleMOiVPEQTePN2rSDJcL3YRnSUEi
1adQF89I+t4RkdTZVyx9kCeSwfA4VWTIw925hsOc9bTwcOsGHnepEJY1Jw+uOqQZ
7RjmH5AUUPLlhjnTCmUBS2QLUmeruhqOWXGi1m5OXsjCmhAgQYNTbvJYVOVkzfsc
KONMoc6kWmUFS1Ayfm3kfcJkdGc6NWURtRpCHdBcy15NvL8fWnaegC9Q/pQmCm2/
e76785Hl6/gmlx5zpbe+9auQQLO/mp1fjNFfFB93J7kd51S/kcGMq78EhNmIK7nZ
QDND6dR3Pc/tq1sbdmWlFliIqpZD8udFUzFwk4eDbxxhxnxnjBPCV9R/xRaJQQ4x
FfWjH99Yeo3CV1O/r7aH6rzB6Ye9xb38sfScCp2qmhQVFOwAiphLnE6V2532J89z
Uw+ZfPUpmPMYqGUOkOM9xpB3U8bQ0dTg0Th1n5+fKg8bgmiKoA45ZzJjbLEhZgNe
XpwXx/OB+0FTb016nNXdoLwaKuPzaiTIXIqGC5tmB3BFgxPM3Qs4WfPS3uqK+rZx
Vv6wkB3Tlhr6oDZTWbnQFn6RUnhQ/EAd9sDR1AGyhwnuQHnr9sMtS+5jFpf+Tydv
vc0IonXamVwwo78ph/LJwi/nayStZIqMHq0mXXtPFxGPBsLd1G2ErM2EIn7o1UOT
BvTTrpZC3CqOSBSBzR4/SpIx/3/yaz2qog/iMBRBvCnRvV6/4fR6RiDFkkJHI0Rf
dz53vnRDvZ7c3EVV1jvt3Zk8BJ/YHP7nB25hGXl/xfIcKfuQr0ZPFqERjumhUP8w
x16Fiy7UuM1fgVqFAxNXhjnvwoucDCfMa6SnU6hC3Lrh8+R0+G0VTYAYq1vNkgoj
Fwfe8rapt3cpG6x0tSa716Plkmdx7smCrXtHgpFhWkeS5trYmaSZ/NrBGO1etw22
k+GCEaH5rMkyxbtfufr6xo4YLeXs8WzY+/ouwD8Kaigk9ofeyFAxGsupGhpu9uUA
pN/O9r4HcLMSU5SuI54u2obrhu3U4T2zRkPL7A6Dym/LYBjmNnbYNTqoNxU9g/lx
Y3wSkMjeoUem2pJQMxuSHEXn+OxyXE8xy8pCNGbJlCas1zo/iOqFYMxL1xjAeEME
MWpfKyZgDN1A25bBZUrEmlwOoDVL1Qyevb5TyuvdfgeVeaq9Ot110Of54a6VC5et
k5cdVwdShR5t1AP03JRaAzJfVyecl0KzRZSfFFCcJh4T5Kle1uD/xv+jZSObzhAm
DeftAHxyzyHSD9Q2g250qlcdurfDxjcKbT+7Ea+Vs3IdKE2pvO+W+5FfK73/rKGI
i3ZVP4+ov8+AimVSxw8PV/mTK1G8hIRwlH+kRw7KZlvvXzq/R6mA/IvW/UgNX+LD
i0ojrqATCoLcA7Y4IW2NvxAIRbtSUfu3sVH9QyL3AYXnj2d8coZJeLv3hPYawlyD
L8WY3fiWYFqBOmc2Q5nmFytv0qB6t9i40hRXgXMLvggrOC0uUEXVdb3toejDnNtg
lApyHeot8epVlzEJiFvUkQtn9DbGnLl4Z5tu3vCxOOlBozIyKs67uDcmPEzB+3zA
xDl86mdbz8K5MKyQ0ja5QFinnKCiirno2la87es9HA15V3HZ9m3h75R83EcUvpNm
H+HUcgOieyMs85F3tekwuWSUnGN8uiQQnsOFFbJV65Z9ZmfqF08c79Ah1+wdgiED
Z0cJ4WFcO7a+FZ2R5CxWGmnKBgzR+ClmGzpdUAOCGvYlJ3fZWNjB/cETs6I2eISz
rEBsVu/1L9lC8Qe6COsx84nlWqwCp3Hfl71ktjumhGWfhlUydyToO1hgE32rzTUg
5jg3vwEPl4iqUtcW+uSSmKNHW3TBi6PBmOSImqu/9VA8A1lWeM9Pi5i1X5h5+YzY
fpAHcHp9UjawpDHCNTIm90U9j7DX9UouV7qtvUiXhFlcTzhG81TRf3tgGHCO5WHq
iztDl9HP3bliIFdVXEmfF3VZBQBmuo2/L/8zdyuRtRtnXZvzY+gzIG7aIGYiAoZf
1xp52ygoo/CgCwjlrjz5K6ldvopZupQUbDOGNPpDXa75IJwNSC9JA/InD/soM2l1
BIES6bfIiqbcHJUVJFSz+K6LQ8gHPauhDQ9bJ1UcflCSAmBqvEveaqLayHNLAuLC
U5VFhvfoKEpLXid0q4Rc+aKbErK2l6Ey3oF5qQ8+BY/KCJoKjMaHZwX1D8D/qE4Q
IP3H6p9uminsFO+G/1woK1ZoI2M2+ixIjZ9NQSrm2+AJ+DF31GqQ6r+myv3JYQpu
jLPgRuECUvGl5tKvtxHs3sOnNtS5ad8UTV9RhNJI6YY5CrMx7fbrowQcJvn4bT7N
ODvmKEKRCibdS6xi7F6sXPvXJWGWm7PVn2puI2Rwf+p/HC0kj9b/1c9xEGXGHuA9
CYoNmvW5SosX9rNmHDSphfSgu/sW684W4Ma3PLLtHHklm1yxwAERli+bhporB3u2
kELTeCHjWgx+N6P/x81PfZ6LLMemS3hF2AjlORoy86HrkRFJnNl7fqb/FoPe9b93
6eHObN1jkoPVeqlLumqxL5IsPub/cNyxc0rR0goMWQQrt04BnviB8QKQ+Fh8NqHQ
ornT+huWirPSFAb9XiPYXgnsOXYaBZvZ3rs4mv85rXifG3WZLP2HmxTH8TyTAOu3
br8BzByOaJ6dUU9qiI5NB7aIyjRC9UvPTK3nFR+hSYJ6jUN+TpkaiXfKlWEKXx46
o37W22rs60kWVntbOsFlp/IAlOqjblJryIX4TwV/H2YBGyF8s98tA2ic3TJs/RAt
dUtjdyQb5JvnI/4Ph+sTk+l+jJc3A5BSbd5Kvd53u660TMJhyuEeu5X2SqU36ocm
GthhLZPXCVb67jVj1LftCMxVoJgYF2vT1E0E0sjg3x7viN6lPv7Hbz0ukc6bGzEB
qljR1q2g7ygkU4d6Rbov6SQSOllr66gzUpm6hIZxyKD0MzCerJfpTqVdFOswvHRw
fJnJF4vEQ6iW+9NplE3NsXRPWsPK4ZqfwHgf7LGgFBfnCMflORIXp+Eu49OwZsic
oJizsT7fv9YURAuBmlJWE5cT2wFqJIOTwmQvxf5LrI/0WtX+I03BAaVqSRJVgEZP
9TmYwT5BMKe7rD428ZK6YcMhc+BCRYjtf7wPxO0k7YNzgfuX1dzAbRHu5h5Ga9vX
JkRaa2BlswB/Gb5h+bes8hTTsgDpDiscD6blgsZU/JfMiEQcfusBFkKAvQOeGNAV
HhFBlWNZraSELfrJTLs6BIIaW1BA5KLIIEoi8B9VmYWRckhQTiaA0ieQsdJ3XWvQ
phyt7pZn/3C8ucllbx0BNAsCWURYV6iuzSipzpHQ5qe+GIBU85991Y7FP1o2D1Ay
DzOcqjssSG0dGReP+Sx5hX2exGg50m5nToQGD7fpl/fhf8nZuNwbUi/fGLlLPSUj
q9oDR2GXi1UHH9+QfODtZ/ZHwEYTTSUWLplJBRTM0ENhxuJ/HOZHJhzHumAIrghp
nb9rm0BeFYcsvoqsBogMwxmON8kKIoLnfOnk3KKGdg2+FtZD1uMJ3X/5jlktqk+p
4Z27DBu7jtUelVQZ6jl/xu6xoGccKRZx2GlNRZK2cAQ4Vbw24aIEjRe979iOGMKN
qT28fQNLYT9brkR2cSnuxM4TutcRHE2D4puf3ZdpXCXYNFCOX5i3uvir7jIiqdYt
IQQwNW/wfTWvZzy7kxuKiVu0paJEaSAFDdRB9DrVLj3Wb/O7qVJCDDKYO6o9+Q0a
4g6wBxdRxSdysLmzgSpgYOctH+FQwFhyH9BEkxkdzt2Uw20GPiKREo2H0wNuVEvF
+dPjCa61IXrgeFBrymeoRU4WB4yjy/fb9EC/RwYQRNqVFXHs9lAMcMF39nfr6MSJ
pgpapQaAArXvn6wVROIA5hAWVte3PFyZlCvyudItyDw6rxU0I5nnl1ZXPksmDCkQ
zV9gqPZZEo1AQdAyW2D4xb3qEBEReJLa79f8FcWkgVlHW1LRORMakG3vUq2NWwmG
dMgpr5kCajZUyu5Yh9++F/ewt2H/NznGC55f++x+1OOhRUiBoI/OX3GKT6QWhwnn
aWLi1VCYK6uElnNKAD97tMnKaaihFwS8q2qUB3dcNqu9DaqePCa2+xE9EdrjAxcX
0IWapYyOV8W3ksRDri59C/Nvs2X1rFVho+NGnOpepJKrc9Qjpur/8Ty6LEOQ59lG
dQXa1NWt20/hbMegB3Mfv8JIwcvbMSnusgtntXCmG+vr4KNRBUdYd59fKrPUmVtN
1AqRJ+iHdvf+dPyi4TRfW8R+vMfa6p8mhg9WTQt30amEVmn+xq3DXfMkmUOQWn2L
BRKi+k0gAEWDypf2ee8iRVRJQioBWrs8Ev5EEfSoF5cJdJF+xfwx4BQs/Wz7LvkI
+nzFOtY3vSGsdstSKFUKztQ4+CQpycR4MQaZ8FJDFYoJM9+zBBPRKjR5jNObfM+k
WqzgO+I/O4DS+q0B4WBDieDzKLoZmpJcloNVk5/nUdyVH7y6W0GdmSufU70G5oYK
ye7GoqdxGOczB+MrV6diSzApa8p+Ly23yb0Hi4YLDR0XO8Xgp5hCi6GGOHr8f6vn
izs8Tg1CJdiNDC3ao38EZjtKuO/srkomG7TU0gJzuEQ9ZMZfWDj0EkoSBWtYl1XO
pesw2MrDRlLcgYlYXnCyONB7Poy9nUP6yjcuy07hLMGLRqkescxyqPDrLYxW8fs5
UQv3VzH23vN0kOuv5cBhTQgI9whu5Tg2deHSSFwT5QHSJd7VfSypffC+S33FE7cf
xby0nit0armtvJ1weIwXXfVSZRfX7o07L5TsIDClt5yWvXj5VM/qvb3XYSUfx/nr
VzHC3ENQ+5kUboISNZQJ5G96K0r9n6m5QPv4kkML+IKt+RPkyM4wPUESmPJlp1TJ
PsRPupsYIuha8CYlaad9BrZky8lJRte9SyG7cjsojw9vy3tlQR9e/Genk5aWRNEm
u7lZHhBDvC6IEQqTISpZZ7AeuZ/sXv/eR14sbl688cLsyfksc8xs2ilDB2JKEGR5
8DcsL4ZF5UeufyiIpjXHVgSlNHacNtBPm53JM5tjsGk3TfxPchtJeG6iLyTHIf4Z
9HJPQPLLiud3Gxnb58CQzrLSfPGvYI86aafNqlV05SOmAEbMPhdqPcj/GbUaET5f
SHzWDBCbDTFO2+OeuUv+1Q9vlhGLb1hb4bEKzS8yZ9M5rAqqtTMHJUCtEiJplcB1
IdLiXNX9X3CTbD31fGRpaSVC6nv2tUgWomUfQAPdO5IKsfB4SUMHiCLoQ7F6IOrK
T8zXtsAVaMIzKK1gzxQJQYQepc35sdtp7G0raI8RSG3kd0Aml+qeqnR/T7/qPgNl
edH5OawGfDelNCxNtbRdP7WwZb0gcu9k0lRVjfsrN9XCQlM7O5LCeH7lCUSKImCX
MSD3SsBHEgNeNw+oixOXw0I73qflBjjqJ6V1iL2JoBMi1+hqBzgijBIeViS8YP6/
tWDq/hEHBuH/pKw+ZmoZbCLLM21PV2JNfihuxgl59Jrs5tBklRpqvx/KrE3W4PxG
d15tbB0WAQh6P/4xYUDypPdM6wzK2b1ogQQdy6h8zvzVuXRBLP0vKJlxA3skJHsr
sIwcyGZhfNCkZGe2tKyQ2SPo6DI6kyDNb6tGOo0uywF5JMUAxGOMmphMnDYWP3Xp
zBbmjd7IrDuZQh5D9EjXkDRykJmiDEmQUFxaC994zxjGyDdzg01acaFbdU1BEo5c
Lx0bSknmVC8b0XIUGG5hRjOkhG5RVeoOyzGvOyWNvlSNPRY0R1JYejrU1Zi5M/Sb
VRJzkdrjbuIVrX1GBvLwMIYvond2XUpCRX8+4CP/9yLkOBRWkYy0nKqM8YlsMso2
R9xrB4hlcESdlWcRByFYkBJH6UTOVgcIbgfdFyv6zrlq6IxUCIPASQcSXVEADN4R
zT66ezXG5pTAERbM4fiyE8EIbI+X0Sd2dCyM51MT1Q9TsMCMxjmTrNB3JQvooiMX
BJWmOYlSNWC4GyqaRMKyNqQoZPrWBzzEZj8ino0YJpPZkqCYGfDBbe9/0ugjqWxc
595gfmeo3o/BkPY6Udr4mwlz6ftmFUMXoTZQiat1hEdQnWwfldct2zQ49lyu5KBb
Zf6ouxzMhS6NhN+8FaugJAbQiZrhuXf0rdjeScD4LRzonHDrAIcBvImorMaDaoiO
aFr5b9AvkQf0z2JD1kKLCteQ8QEYxJfhULbcLcqRUoZLqzwv/24qyXecpkLWtLIa
uRUgt5eERxLWNeheIHKakjMEVHCEVr3imBMK0bjKv9e3HwGPRWfulOz6jm+28VKK
jYnW+Q9/iAdB6oDrVo34dUgtKANMz+XHcUKzQiuwfpzaPBtPFMJfdEJ3eRvJZEDo
ZfxyzOltoTV4Os4Gx4l3s3HPahRXzIZfocpEOuRxcg2yBZ5wEzEzRVgmMkID0toF
FMd+NhiQl7CmMnv10TrZMNQJCCfENTkDhoErZx3AGg9TjGUm3kFjEWO14OVEnFFd
1ICgb+QL6FF71KR0eqo1mTmJf7CX55+LEqM+9FYuUTtqxEcS45FyzEm+Vgslqot9
+M+UsW3/mS90TsFRxJ+V4wqDxMTI3/S74n3iYp/k6gM6cGo+ORj5OdpXwqgJa3LX
MNGc49rv1LbVJ6UZ9CquMU2TjrTNWiIdgA0WI4x01Ctg8RRpEmoyJG61VIjWUS+o
RLjRNsNF1SSBWyjEZ44qke9rkV1qvLklL4huvFHDp+Uf7fSUR3Jx/JLH6NxmERMo
MBr1Q7Qdf5+cKaRJRcPApN3RYwb8dbQMzuCSuwu+NUAPqFmgn1mOyTiRb0zcAcOb
Wf8P/WuKzZMJ6z9Smc5fwCIi4cwQ5bys3I3dZ3RJnqvkJhzcqyU/HZYKkY4o6uHu
IjEzuZ3sdE2duuE8bDo8zkWQkyIvpBIyLJiEmqVNvECuY47QyGkQIz+SERgpLKeh
e1b1yM/+otU1NTrf50dAEn8nonFsWcREeBeG2Dy0ZY90jbCcd3Avg7/9bQWvPzis
PxviFPPtm8Zz8WY7pDdt1QR5dnkmpuym0geZzteTLZGvzpPsGNb+3s5RJlvyHSmQ
V3x+reP4GcOcdpOsjbyZ0NEeESIicmpzfPe/iKrG5o/3Uci6gm9t3u60in1OAwmJ
sw09XpZdTLzFMq8P94105uGZxZF5+hvgLKtMm/nkGOcgvDcwsHZCEAQb6UK0tqu1
izQ9P+oQVftLGw5MKRrVO4a7sX0L9vB2EwSImMuufiy/yfhexcq6sZyzBip21f20
YUiwA13daurKtoiQZx8B4icw+4XroB1+ywNKQQ44XAsx195nyTvVn4zv7cq71V87
HfRwCM70nEoW/s7MNhPzo93PRcUlWUg2BkHbydV+TvrPYh5V2hJ6nNeAlu0FF9Ff
zrgY5H5s+dG+MGCKn+72Xifq8IzouBYFAdNqlTBm3NavmqVT92t2V6Ape6z9Eia8
mg+ZW1fFNxLWlfpNYRMkL7xWxdjMC4jIa8P4KviIky57Q2ZiuFCoSti+uM5TW+mo
C9x+hVF1LD8Kw5doHh3XIEAULujUZ2ZbJi57SOkVij9iOIPiil6NzoVttmViH1Kk
ZWOHxWts9MxToAVf5yvc9NMhvU7Yg2/DqNSjnNyhA8qmw0g1z+YNBthdChmWP4kY
poUyOLV3JFImy3jkGlNyKt6U0CpWi5dep0V48IGCuJOfCJZ3v/PXSjRe0nkBQZbe
bvtrfG/jEQz8L1woGwQkaX5OygyOHbha9faNiPtxS2UTwSj28FEXP6TOxzY4AifU
RfFsgky7zFU65Z1LWrxHsiHaHSzy/ZZur7nM6DjwPh4bLJiufSzGp8WMvrj0Byo/
W7noN5rq3M5wSqrItfHXkkzG3v481LiG9Fdp4l/OaHPbcNmCkVEx6Zix/UXRwiUW
4PZKJWqp6CsJJ5h87I66C9hPlSeZQqTlqZQ6YyjP0gDLZzYsqUGQ/z/bhCXB4Pa5
XPuQbmLIHE2GTMvN3U7YouwDhlyPMyu/9H6lVwziqYctUuea8S2wgp0E6W04QFpZ
QhY9nXMJpOSCcBuZCB4IUXVDXnqq6KyH8JsQjmXKaRp/pHwhZ1RgwokvJjxlacAZ
b3WX1IJrDtd/hi7vMd85QQ5vkd8pkERaXou8CJGUCf/wdQCSblHlYIFzyRFupHq1
A8qSmqdFAWCpXgTOGTZv0rFUmcB2ZFVtgpIApufjgU0ZvBvR6RVnflD5B8GAYJqp
6AoUrCmIZrtHVpTH6fO/1jUzWrU6+4hGMLsJPZYOIE7ovJo9oqIxVXIs93UN99Ca
UYZh19BgzQDByQfbYZ3FN6Fp/yb5XmGw03sKEIpJSii2Aj+FEqG3wuHOv9RoMLQ5
a4NiEp626Ht3O6Lgf+tf/8DT43JtY98nXLuHXdgZf2y2JAEgdRdrbaFN0JxoWjLU
+vBea4890nmr7ih2kCBlbcHtQCy4DLo9c0FWMZ/l3InOhy7AXQpPq4ZGe/OFapiO
5aFeXU/zT3AE2u9/y9wON3oyebzGkTsrORhh4IF+BRaF8nkDVySdLdNptt8GYusX
4kHH0ub2Yks3Wnwb9YHdD2vO83H8FzTXLXFkvYLkK/eBSC7cdq2ocoWdDAn1+R7t
seQNt3iIjsAL86DZpF367nHsbLDJrum0IfW20ejX/l0axgSoTBlRio133hc5m1DB
MYQxluSfeTtM47vmGvpRrStu5ijw6d8FF36AWmm8I/kOwL4FC80hUlFujFUcdKze
iAAEgrSK4TAD5LWRzvH4dZlYJFanPkFf+v7fnH5qKX0gvOK2DlGN6kVuraUIwznN
aJhd1Ahit8yvFa+y4J8Cd4O/20ioITrMu/VCVmLSkuNSJ6RH22KtdXwRQS++Q/5k
Hl5LjiRYz+qVLQW4UhGxrdIHtAXoMClnVyC81SxywgGWWqjPy7k7BL3oWnAHWpFy
DArcdBOJVY21iN63nheZ2P7AmvgaUH9vLuq5JKFWnRM/LjN/xPNItSn4DtIrzh6R
X6IRjUNuh2raFecD0YTCczOM01rW8N/Jbth7V3er6wJwZ0eDo/Xgg7TGdmPD3uAI
kxqpeZXbp7a1GwrTYCADEGex6gBKWeAjB/HDqPEFuR4wKpzm9ukhEMK0+VcRZ4Em
fXHqBxP0bSm9+lwQoOvf457Gf9GhA2lCvOpxLWEFBTS+OvvfO1eD+HX2XUOchC8n
s89OoG44Jstdx8LP7vS94/8fMpk/s7fekK8rXVMdiCW1SQ2Fk6e8kapUoIeR/w3R
vtucvfI1swl7S6ufOc1TQTl68w5Ay3PQixgas/RcGQyojbhu+GdvZXK7A/D1rrbo
imXGA1/go0k9+e7muX7UhfOh5Dslq1tk8u7ATb1FnEGo6OqkQHlEirswQvcGIH0r
8Q6gqlYZG85odz0Ku3OCIzqOS7KDKth4oYGCSADvXBEIWJRV9hqokfq+LxsUKEN9
mgQJj8hevHN/M/HfSUgjXgtzQbiC9LaNA8Tok/GbyjDyH+2XAEuM+xRK42aFLwip
ovMG6nxvd1PZ5nlNJWbNJvSgHnsOJZF8V+QmWIurY1MkfqnixY6m4jIA3wFYtnqR
U/V9gInVcLraLl+ILdTaW/xq3D8LVKZAOYZ+g/VekK8iRCYd5JbaGgrIapEE/9bI
t6I8dm7kKd/HRPT7qXQBzSBQ5b2a7Fl7kGLiihZSBcXYQ7xAaFHPJxdgRSgPmsmu
1w9clR+Gg9Wcv6+kdgF37IlCU0U0f/ediC7ZJx5V004larRuslo/fhzyykUi4wsn
kCOjvVfFeNO8H+kU/Sh41d9zRLUNkcBzNjKSgWYq+cgCCAD9aPw7S91m74HlJt04
hiz6LsWBOMvJhPd6F1ZQzx9VQw9+2dNx8KttLFv+v+rDoYFSb81NltNW2ar7sL8S
bYSsXA4qe0WK1ycvM538dQ4RDav81WFw/TheP50vVchIEkQh925gn4zACvxCqAXh
LANX+20FooekKKsnP4T6T7Z1iK0yD7vU84mEAhKQsHM7bFIDDCw/bS2ebTu3Zq60
yWt16MPKBEbV+DQUYL2tc70P4eSiU1NN2saRbttuwZJkTRR1u6tq8YqQ8F5be/Fv
p23YVtM+0iXKMYDnx7vS/WqdHJFqWCu7Ma0H043igD0tARAC94FsQRC0r9rmXonR
LCimHSdVgUX5yvyiqPbBbw==
//pragma protect end_data_block
//pragma protect digest_block
86j2l9kMFAEKBnjlMuFcOKmJJXY=
//pragma protect end_digest_block
//pragma protect end_protected
