//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5J1NyUeybvNVfF05F8hk6LLSwgXsWAh6z4F8IkHMGAPueTeCFzp7VS1N1SljGZuF
3GQu4MTTBvN7NGsCuyvZaYwmS8vZPvKB/Z9rRgCiKYkU66ZIWUJgXMudSfqSBknP
6cFxgO0+igiHPVFSS+EU/ZbCqHIDRqY5wniigSsSrTUyDb29Xs80tA==
//pragma protect end_key_block
//pragma protect digest_block
NwIX+0hrMEAmJn5IsF1l6rRlAbw=
//pragma protect end_digest_block
//pragma protect data_block
O1R1piwdMRykfEPvsTf/JaQpOGkRW6J90eSjiwAGASj8rV4m9ahgr+U1BVNAgCih
taECy8+l/4dSc0XzYE+cTUzq6DbvTCJSx0xm8uaBdbAiK0Kf0tEgRZ49FsZ4ewat
SK90N3Akb22Kia8LIH3/gSF0DX+EkE5lWRfAIQ7i6Ui4d60YbzFWgdDYsS/qKb5n
6bIZCzKG6N8/G5fnScQE3Iuqv4mrdXqxfuKaRQEnVyoVjdCnbcsJXPgYn802s4Ga
SdslD63i+68LFklzwMMLW0MfQHvF5ROQZaouvUxBDTqLIBcjQQjGavcVTDDexMPT
fRDyfMxQLaismhTmTYwaW8ASURYL1kdshwwbFI8MidLlBZA0RkB4Uw56790MXmc8
WNT5uGeFzh/8qguOURPOjKjQvbOFNDf+9MJ1rfK8/M8Qbz+eoWdvU+8lBdu5bkH1
RgySx7SVo1DR8yWDIEsmPMa6aAsbk8UzVJH8VZ51OxpcMgPXRYxgwoOZ5041Ewmn
xPuK4rWOdhKPz9+DPJiydig6TH26VLEYPBtSdoD2shQP2AUfl4YXDgt3DSCkd9qg
QwGE48FxslXPhuchJ9jRlquDqkWm1eY/Fa6l/FTOquTpmURL9AeVB8FtctuECoNF
FB780UzxxEOM9dwZPQXs7JGxuPqv8ZFu0CqlfkcI20tFhuFhukur+CJqW4huzSnD
kg37i9V0pRbiXVbJqJPWl4tI6FyjLhpdvLA15br1+JlCZeM9C6g1ZhtM3jtQ1QxC
nRErS0uG8kJp7puBVS6Nmf81VhroWQoHdbzR+ZyNz2/bgwyXQr71F6wFuoJUXzqJ
UAWSQv6J2+s3XCWYARtkfYwO0Zn6zWI+b9Pd85EaR8hLUjVbwXb3HF4dPTXbP/Kw
8D1/7wpv+xLo1ACvJ1SUssDw5W85GfzXjnx/PDazTgVA+UkEl4n1spcGjkMChk3G
euRllHSRo3bxapqVWZhL2rDXomZqSeIDN1xSp12rt49AR8SrKx/wjlth/hs02W29
g63i/IT5T6LCQUVgy8EwULf1ci9IMnf98chKGO2DoBHgrOyI3tr0Vf0dgBaXNfs/
nkDCqh1HRD4LiEEqJL5KVzloj0EdmsrriPZu0tJH31BXk1uRrLAV27KwFypS5vA9
7WLix/3/evBEYMOomUqTruNKR/X46dAzi0V8UV9OQfDr7AhgkcdgMYUzcvisOWP2
o9Q4TdvWkCZeYFhrtvGZMGlBO14cLlM51dxKdKYkpnIdddKL8fMkfne/yXn6xnf0
K6FsfygRpDf2O7FhwmMG+j6XJBs8c05Wdo3SnvdxHZZEHNxtZ7aSUjHW5ey8eFxV
pyRYa6ruIqVgDxCoRYgbcBuma5u2zNPzwiH33zCoFyPtzNXaL8RWxEJEcSOzmXib
/VlDHaSfH+E84KKww3fOunxOoLI7MQeAC/AtHBfsFFXvwI5IeCk96cdT7M8HGzNw
mHiiaI5MVV3jLiN9K4MTu3unKE+VCVmTkHSu9oqRGBgxUaIrly+5KCrRWTT+yVtO
Vd7yHkZFjpw+3H5+Yt2l0614f9lpeMb4gLt4b9C6XK3zSxojv5FXCGz/wgIdTpI1
L3nyz0jZ5nog2gDW+oXerSxIwjBIIzFJJqnPRgWkF77lcXbwVdmc0sBLa1FmXc17
UzdXhivv3meS1aizB+50k/5w1uMyFv0UfhdIg2zRzWrM8GmY48N0B57CEvB1XYyz
1Lq6QAarWhGqOai8st3u+Py1XdbxmqmpcikNU/+nCYTznSyuj3+dwWKJXNeVD9JR
JkmQTSo8bvORo9LM4F8fUqBV6yBJqhelaXvuvpGVIEqWWHwL44sV1xX1u9oUNPyq
6Gk1W7uTf6sjO8yvuZgc5TuyyH2LsaLToULRP3PDlL9c/v64ImCk522KwDWlKEKs
wx/hfwluXvcle6lR+iZEakPPt1A7YxEGRNN0yM8bM7gT8e1PWfzvYukUWj0NcNJt
6SV3eiqVhP3Rq10ztNwpnwC5AgO3t3vM2TjmPnEKK3FxGSzhicEvCe7OOtgV6wn/
ObCMt5gu2Nr6lgx13mUxlJHEmTtJitY6sfzOVMbHyCRIyyfNxzF5CqfP93viKdLz
VGiTNB+iv+LH9SNGE4w11jOJNnhKBERaMhpjzBR1IgtHd9aPyAXiz3ElJGWYSR40
Yfxj/DItwrOu9KaphSyeoXr76e0PqARt63n/aKKKnZAnBl5ZMSYiLieZRKHhEq5c
pg3Gsat5XuXTLVjFNeSuVb76K1YaRvFgQ080EsM+eo8n2n1QImW3V5pmZqSTrfSk
/mG8TwrrZUdeI8hFGQJWegqbM0gKMr46ZbRR9P6w5AlBiOfs1SskhcR7ic0IfrZ2
GtmwwQG34XdD4ziYuxsRPdNGoT6pj5nAnlyvbqbR3SuIbBypgFO4LZ22CtiW8+kO
JxvcNMvI+PEOQGrvSQ5wWKhiwZEToH/h5x9ToqhfhD/U/Yxx7icHSacM784jxMRl
8ACqSWqJfyq/bt9WOWMhk5wTzDl08HKWYMj+I9Xf3wbugI7J1oMaCTAQ0dAr5ScY
yKicmq2IVjXmS8q10PLGjTBjYl4wMXclfx/OCxJIKBLW8Xabg1HfY677BqHsk4Y4
Ci42K4yItJljUvaiL4vX+puNmE7DW3O+SbozEVQd25xQcp2H8UkAoTTA0E07LoFS
1h7IUHVdsnbS5W6lgZiQ3FaVscqPCMB16ypxZ2nMrNd0FsUUD2tPSgWVXRB3DKNw
v7X13Z/ufs9vZoZQTbCdhLurWBlqM2wixxcQJpuWT8m1q/YYEMDziXn9VpJXXoz3
F6/0h1z9MIU8VddbApeg/vAF6jHOCIJ13SVI5ary5jbmgY44B6RFxH5Z3T4J7e5F
6A6mZ0F4XdzKR+zxAOdlbpRdtPSUlZaeAdqYoM4lKvy5DvAmHmy1tFMoR+RuURPv
Aqes6yUHArvwwBc0PDCC5EwLvH8dSL6Hchc8HXdnaJPcvFLvZKxRgslM5FByaAtj
+igeho7/mofKHNpxTcSzWpSO4gzvtBLgXF+BUwGkZcvhzC69H6RqGudIfWAMQjDm
pGHjawTZFXuCmYrH+I74OqMBAl3nyq2UppzgLt/uLnqO2NpMXaUVYKA/rUFuFoSu
gpEFlw0YFDItxKSIZvude7uB2a2E1P8fVBlfMOvlYI7BAE1qvwjous0P18qNAhsg
8cyj+u7Rz2IiftfTLKfjvIGN43giTtE6ba9S4P3eaC2wdcasr5fJuDKStmXj2Cxt
R5F5+ZFN05lxWSPvrhWRieLUfFEio1kltl88iteaNLxXgqol+h2DOAAm43Ew7b8g
M2EadSKZAqByBIWho/PAepjlR0JoTELChzOw+XttLfa5KbbknJOTZlv1oYSJWPqP
rYdrFRIl2i4L74h/Jr23PamS1RXhrGSYxtU2ApBmUwLu/JeD/hmKXc8shxZSRzPb
dokzHyht1RDJAF5Or+TcRsvLMzX4Ii3MnLkyg4Six5wvlno9bnGkMVb05K3ODIPy
2zLNTP0nEx/17dvQ79GjWZ2aO5VPMSe2F7bfY2OhE6nLR8QhObDhXmi1TIAv1oGS
U9gKi9ySs9/IUZYFhXAYtn+txlwwIl29vi3SAazV9n/B3zqJdFP9XZFa4dO78FXd
hH6eUuLtY072o0kvv4UzimG3Cb+QBlBiPfQq+13EZ6H5uhhHRaZkyG0niF+augNr
7ggOZMD+GU1ALiJc2CaV/CttkpFxtFmUHIf1lMr0/mHH9O6ACOXWi1opX4na/e6A
Hdcn4ML9mjphOQJ4hKq38RjPMfssqGFzKGM5Rpai2Eyk4N30gcd/jpA9mx97xW3Q
ZXnw82xIECAigaPN3leB0GCYERMYcblwOlO5NlChvX9E/s9R5VnQCBEbaRkNs/4y
z/eONWfpBWdByNkbLgjjzhxTyA5Dba3Bl9PTRmN24V+LsXGiuVIMNFxi2bOXywho
ru1z8q/BndAKxQiI0AC4WjKeVE8kEe9PHZEWuhfNG3ltd09c/KAJV/rudw1MgFpD
VVfud1OlPQYRo1c6qi6yN7n+dyWxxZPqo+84/CPY1ho379SMUZOpwzTgx4oy+Vwg
ZDArjeQ1jVrk+xTa4i3XmP7rcgzaUmfl0BShQ52M818KSc7EnylgtYOG+WhZMqXI
lR3COHhEQmxZooC0H8i3nrhM0GQm1HYxhe4pN0506icDyJU/1vfbR0l213PYHk0r
Hsh0x9VYzWkrmtY27WidhUGqscNcIDk+AA0tzVLKumw7A4g1sYmhCnrQHHQWwGsU
qfrRRi/YbpymwwR4/laBMhleiXIoLnn6NqWxLwaTrQTcST7iDfVYWj4KQawBytaC
z0RvwT7UrpFUVpeonTQCBIBMrJMFPiOokwuOT2DUaG9zLtldtU5+854VfYmfj63Q
Nmqj1UupJPpZGmGh3EBhiL1S67xtVhKPkMjKkyGus2DvSYrT09sBbiS2hrW7TZ+h
gzlff0sMhAd+52wp9ZjeCXUXWiDFGQbdS8v7cUh4m619j3k6vFDVtO9OR/pWxe46
YwXbqj52Gy1Uor35MeFBNRk6Phk0YH+taAdTAcRsbpBCT8Md9VwQFbQx29RleHJX
1GRHagcgWQaJ/W40juSmaIWNXL0rdXpyvFuV4QgslzPGTIwSDvglYH4t4FFAaH4s
QjyXo1Ycw+0UNwaOW/iG3tBVZvczhDK6e70QCiLUaMJsGA+nyykVTi8VwX9UlDBC
ZJn2I5M3AIVnCCpCifGgMKBOEYWAAJik+IdinI5+nUXkGs7MAMjLlpYE+S3oOqDK
bFSMfV+m+Zgkkrx7PxIduIGype1k7hPacqmLLJA4BH6ruPBCWA4poGyZbOdYXfxW
LGr0VCtEiLg3Bvbr06EopZgnaUBnsH/uBR0WrZEbXis5g13gRWmdqrmu8kN37pzc
sznIavtdAHsNBepnbCgn4ubiFKt9M3ZEVmB55cfGdGKYhsO6ElkPkZVGb/wPHZJf
jUMOwtXefZLcLT6PDW1eqQUzx62ld8zyxBg/GeplbvFBGcJEoWX0WurFRrM87ONw
KNWNfyAeav/iHCPGPGyX+HHBP7lXjNmvV4iNayoAb8PEUoQPqiVQxuMSUd901QlX
WtTdNVfntrgKcybh/zAPKCQ08g9blHjhzUyCPMW1SnLwHNRlnxj1QKD/FsVXMKUG
KHLDf4tICHk8Y74Gfcc2gGe1Y/rXxWwQvVl7fAtpIdd4xJ1qFuEZ5WMFP8APJre8
VLKkqlqE3dPkLQ9sE04LzEgyUujyCvt7L65vtfECTot6TIWlqAsAieU6Sa2PRnSp
2YU5zt08xBstQNsEqjybO89b1CwbyyIMPCEnmp60/pPi1Pvsf0yrGpXKuKee1EfA
KT4yE3lB4ppxSM5PNyNGXZJvVWZ6RQthGE2d8MNJoAKcDEIRgo6ufp1XOzvtIldr
CJTBZiU0GbIvy/gR0DIdsySAfaCazVn4CZMbRiGMStnrOqzJ4Dwm84mWPQi/hIbJ
WlkfmEv6z1Evv2DpF2ztQjAvPPYNS3k5byqjHhsbzvSMJWIXCKq019LTWnoK9DZL
Gp2jYHBg/J3jnvqAA0wES2r1wxQAOO22SvEDi3Gs2icPjSQaRbff59ndxLK89pQv
naecuebUyDN9PTwkcGwwhCZ1OHy4G6+V4r3BhcDZJtKF3JyKb+yuU0EfA3/xJzBJ
ZLaARvzpgN+WA0tioxzkbwwQwINy7sfc+nsJsxCBY/M6VlMp75I9T3tNPK2ukL6V
dg9m5zm5XTHgNgXS0RAahwGBPBaWRb8CpxpII9JbWkJIXyELm6e/D/5tOiUd/1PR
GRrMOD+LBSocIAva7Sp1/CjjL9KGpdIvihb98TnNYmNSzrmI7eN8n8WFKZo91b8A
czNN28OsrFC0wyp2HLggJa7ZHzB6zpPYBDzWshsjayH5Yp4z+S1nyG7gSdzmy08i
kdWHznBB8hO2RRqY6VLgIFVyKPMeymxLFzyWrEQw2wKRW4wjgHIIWNG0zSNKG3ub
L/pGa+PyF6wbrWbn5Ttw09iSfJu1vHZbsyI4P9nuD7bBzzubS8YhjN4QLEjYFDHu
v65zMgZcZ73BV3jJm1KUoe06a3WJZCxJYcPiPc6WSAKnbVULqO6+7aW+xyU0k4T+
SrlTQL4J77OI5XdfvTguu3n0gs/hUw8C8JNROCIjQPhWsJF8195NiVa66yktX91g
ThFT+abM6F+wLd3jilNhs5M5pmDHSykD81eTZtKZcc3v6hbTLNXan+DG6JA35DeV
qbwNoztz3VFY1VMfvzSoZebManRUiDCcFyN7o/0+K2moazJi7QwqBBjgZ5VRLt2U
5PLrqQ3H7ZVDGp+26S5MBQGG5S4KZ3abtEHfx1fRse7Bx5N27rfH6Mwg4cSoU+Lp
OQCq3jSuIxXAOoCfrYNTEMnt3TRuuke0fUXbQUoIYNHAeAgaogGPLjkQ9HDTzCeC
caHeDMsaU8ZQXSfa6IoF4eD4cOWa/Fh30n9XR1oP1KAQKDJb4yDjRnpu9gA41IYu
3IuSjpqOBSFGefQpFp2wCZIeUD0kEGkY61pNqtTMQJkXJ1t2lt5h2WpYfCpJ0usS
SsPtD6Enzj4aXbWRbHIBuCcSSlCSc+SYh9gd3Dyiy4TTORFe+bccHdNYz7PrkU7h
mKy89p0wlRYqkafnxQGayTtXQHEE6+H9p0DXrhodfGxj+/Ustq4Oc0nPSSu2OAxv
HKM5z7AgQHge9EKdyiuURsv+NAONwbEwyKgVt9mbkDemTPvMzgJAMH0ca2FgUxTH
kO73BHwtkPzaPR7MrABowG9ezCQC7qo2No+k8MQdibaKV0NVazgIQS+cSSR6wRLu
uB/lMeMFl2LITmHtj1iJfvT4fBeLGYXqaIJsblgWCcAIu4w3b7Z1P3Ov1nW1jDRh
hCNizezC3dFCxLQJnG6RUyUPrhk0ln+OqIuQvtAoiJiOVA20Vt4MTQRy7HvP9Ajq
lsfL4Eh2VqGaCZo0oe7hcgOT4OLfsOcbZMy30veptMpT2oWcQoW4SLyPxTbglWzk
phG+kfLSW7KfMc/ofprW2gwi5wqYNFZ90Ws8dogkl1zzjsJtK6EAiwYBRkmPWQZc
h2nP/p2Nmzau6hSLMWJpQ6ZSzPTrL/Fzbob6FvyjfrbEHJpVJQggMIxek8EdLIw1
3pCx8WJtVH4Cylf5lVmc5ipBUlNG5P7AZQ01ntXMC+xPXMX8nIm15w5tk+50c46g
u4xe21O+Igw616ft5YbSFKbhqYfOlSFPIAjLggy6Mut0vsG4K1SBh3c0BvXVU9qE
UWWXvej5a+SYFvwOIBfhNXnUwHRqB9PG8x9sAZSIrWXff8SqJjHDieNVsv5rrNaF
/PciGCkw6xm4lf1ZxypO373UZMXcTgEvqWpvyJ9F5Y5nBwhbYJ4IfBbrvbL+gbVS
Y6qbqP8aQ5Di/JevIEzCyPfq4LZhDYb3njXtqSgMI9PXXiZ/9cyRAWTK0dcF2KAR
nkJcEXAhfAWxEmstwTsQPJ30q0Du3QL/q0GlY9m7s2PYoz4Eqtad0Dsx8LIrtI2H
QHq3OU61yM3xllI87g0rXXGDPLbs5K7CARW4KAz0is+6a1QW33i3X3ohqAlYi7uX
tB5rwSSevs6ryhR16t9rOwi9nLtp33qxnlDrUe4TIU2K1jrIp1QvAFDkodyLpE85
PbGGEfJb4PWvkAar7zlDfhFkR8T+gS5Caz1ktMkWHXYAI+sNPlV9YJspnh0ENELa
+WILT2A48iq4lvUP4p9h6zrsx9/kVV6w0mfYlEPyKFq2wLvqmsPEdjUS4MzVrhDm
p63XcMW8wtvPwtWuyiO5lhMX4Wkdu0O6SNUEIRyH5RVeSfuBiae8B8xNh+BGwH6k
gb/0pWwoSr8f+fo5FAVUtMRlscJY/0f3jPXP3cAqIQmWXKwqDe3wVYRyQILgI/l/
u/Nyw2oDYoLPOqRAtqDxsMobIRn/X/mHW3oidkAI3lJfS/fCUufwib4OtYIYC6KE
fm20jhSKtq0+HopcX/1N9jgyUEabwlrPn01apkuHgVK78SfkuUOep2tL4M5KyuyE
4o0riii7Eq0pnjb/CvoKPVgcB7HZPoe4yFNzUSB3FKLUTnGOIOGYDasH2swVuA92
wl1r8oSO6nFRc36oHt7FS1HbOgFo2255APBCpHzunxCOIF8xI4IGN5O/HtNkUn51
LZqSpLAyshqyhr8gL/EzMJ/Y68a9O9bdchAyemZQ6XbVXwbAVZEmW3/MfZp906PO
M44B1kSxWUo+80MCXxqcyc8WC7Fvx9k3X4ZEmS5549ozdqv2jDUPc4WE07jByISE
uO7QqsG51MxXBR6X6Z93+y3h8lzJ4ei62UhJP97Jo+tSB+AlRPFz1z9plvNkkWiN
rgEgK91qLBLWSp7MzfYYfFjkqZIe5R33jNf4qKz8ikPNKLIuc11fb2nYXJ08UhM/
xm4TwaFXpPZYtQOZjpeqKODIiWwSQou68MarEO5KgmXvrh0fKVfqAbYgcuZSlcJc
kPtds/6Ljr+u14M0MqKVgDPlbbRn1rVBzwuxObHaTFwUH0ZghO0kIy2rPWDbqTsN
vw0CJOeL5QGLWRvYSsBH240LTu7TwelARQSO38KMyVqvNnatKm2CSGauDd6nBTZf
TRxEoo4JzTNmqT128szWjSZYwkZ3jqnMwWvCZnHI08K4MBVrqfki0j0GUFs56HzZ
p6X2khLrA+tn/m+4Z+402Uda/8CT4xTrFlB4o5L//LG/W0tLshHbdZ6RTDgrU054
DbeED1gI63DVyldMw6t6h8ENKTbrNeUjlcJR5jVeHTL2QQ9KXxYcJhjV1I/ku/Do
jlXTzb83Y5X4YGFjZeuaGJhLJH/reb96fTA6yCExu1Cl09xU0iSGKuI/fCwNf6tv
ongI2YGHs65rFuAFSR+9qo+AAKmjtc5qzpbn+FBj+H17JlnUqVmOkMIr9Apc8YcA
wuegfaRE5+fRHFCtVo6NtmeI5S9BftYUo405r+Q0XVzNZlf5HBK45XE3JgnrOmLi
4UvXdblJ6Ic1g5BrvqnxkV1GddHxS5unCHvswsQ5ahH7IVwXZfZ25Qh8wPrGRnlW
srGQz65kV9+jgtY/elee4TLZTY+cqsG1DfLI/5ggVbJUN2z2iPDVgVfvfUTPmuO9
ozSuadIJ7M2HCOwOVLC/prkF+soroYlYVlWoVS5pnqP0PKfdaF43uggvmY8e2mbE
PLFTU5q/a3euUmE9Gw4UPp3NNjg0IR2G/71aJl7G8k+ckNJDqt9oeiSTSa5i2MeG
sfBkJs/o81vpctHH1CGjwTvQ2XyzuSdQgTBLoXw3mF5myT8sD3530hhBPf8kE0LC
XZuKrfRv7Ryj+2f/tNp6Y6qAwmLeQoWAVAZ4iJAtBvlzC/9tUC5+QBTvNPCYmNmI
g54voH+YXJds5aUWNW1tvbBHIPJrqykK9bK94dvPKie6i5xqjbv31VfuV4YMteRb
fI+MVanVKP3hgQrMVUZQ43nZBX7xsjFQIpmbomiP+lHoMW2JmmSpgDtl0D6pcf2A
lyu9zigLBwREksod0TSyWL+XjVADNdky/BpS9C0UogE0OqfhxPSvxLDalbwehig3
xCh7r5taC4ZrXkK8gyU83bSsD3HRYkMW0tPqSKx0nNgoEu0XVOxYDF1MrpuSyNsS
sUBGVu4gJXsYmt+5zLnc2yvxwz9h/WI/4X/ikljahDYTilrBTL6zWxHgAwDtgke2
Hg+OmXTjKELmI6UHWIlKvilTVbWRlxZxEM9+4WyZr3iUUxCMkIRcsqkUPcYpjGG3
Y4GGUJqolc1SsNfpTsbDJDJEmDL2XNNf3IhD7cazEoQSCYTIQThoFL2Y1x+ufi59
Y3f/1LigyZanVh9CNFPctG34plu8I1UnS2eUzmCaKbNj7Zbuzg2C9FTpqjw7YmNQ
928qZD/i9pL01yr5Cz03JhNlYtmjIADE0rT/zrXnJTuV/7NWs7VHAo5V7CDIjtPr
V0dukroLofLOIRdHwDlC7z/b9q4eI3vxjSXeNFk+tJ6w4eGyWgOn/LkPHpJ7i/eE
OMpl2Djkl5Zl/yA0toqeLmO+CTsjkaE0dL1OOTSq2jGeq2iIFcALYejAur7GioE6
KFrVAvJY26XemYYnDe0z/tbp/P4J/PqyKAtLms/zpV77pjs7N7PXfA4PwxZPjMrh
VuiSaDkmlapX5NnNaBn05lKt7we61pgxdMpGfrx0mqeAASgSHhaAu/atek+FSPCw
ky1Xlail3Ki73uzmWF6oibpMVpooGG8sqKdLBOgPG5FljnrQpfgEAS59myQQqTo6
+DLFjnp8+2FHEkIvjLLYu7hhDGzidHn7S2mwmMBnXwJ7OWh6eDcB70qM+V8+BcZQ
lwDUvVkJtZGb9G2LyXjTpFNur/mrST/Tt/muEyLmdrFNpP4iTPMUaBOacfbJGict
MPN7mhc/oX8fyvv/x/D+eL2qnKwYr59RXvqJYSb/hcmOCIU65M5cApPliqkHLepX
VVkfzR6p6RhTXip6amzAVTiA3Jf5JI+vtgYXvqQ7Tcy6K0WFLTwMV0KB4SQbyl9w
9KmLRHmZl5Lkwg4ldWczHgjnIktaEzP4OEuuA5ndYbSWtynayw+RwyFj0AccwsRq
Z8hQcmU/897aeRgJBtEpv/a0MnNu7cHP0iwYiFKLeYzbNVF0/vqgsC3EvcRQeQhY
j2bcm33EDb49k1XOJ4DsG2riAisrZAq8zmGWEMi9X66xb9nd9BlFjdmYQsDAmxKC
5PdJ0nuv1yWdeEhXzOPNGXW5J76CDFkj9o003L5gSeQPeM4S3OWhMOD7Ia81H8w0
1au8eZXNMLMTifcY49zjdLbeFSjyAg6DmPTQE5FE+MD/npqxiobrj4BgfOteAAPd
Je/S6mOiqG57n7vSDpk6IpScpu+I4BUcBKWq+rmTNU9NV5mWZjkOzKR2bVEOT/v0
x2gq1FchXdFCBuUNgDTfa4WGwFP2WI7QRABWazutW2DVx2yoZIrIgx30tUJbixAg
+JhTVruKVDW0Bn6fGxkPzrpCIG+cfnZZM8BdzLkIOF3O3yw8CVhrEUcIlZSKoSv3
4GB61fAqRElcFjG+ek81apj6V6A+HhTlPZlijY5pg5Fh8ZVH5o+hMqRFHojwpX1J
1w1RK8bpL9q9LzuuHZqWxNL0agn/yIMFdh7JwgPjFmK27XmNaJq8xZVp3fQqiyuO
aLz3+/iTISFvi2Q2dqnLOPFCr+IcyU1uIR//MIsYTNw/4o88aO+SHVKg4Weu79ww
e7ZXkEMCJWON9VKkeOZFnJORRoimFdhvh2X7pUurb4fLYlSbQcda7w04RyOfBTWu
2qLJBdRb5loEJbPWmc1u6U7xBDqy50btWs278/qF3VwR2fHQmAfHN2+pEWUfVUHr
9+OBPrgf48N7TCZkj4PGpZuG8eYgelmfD1xJQBbgqR0J8vsp1GsXkJ20z+ueoTDD
ayWDfBH0Kgt3ktorV+GAM8cHDlkcpYzdXrWXJuGWwde6Dj7z6AnNLWw750KP1EIX
XSrgF967DDiUx9rMa/aPrK7ieHroN/+eXwIUhL0eMWnlYhmU4uT4eig4/TiqQG/U
poWdHEV9KbgoP+wOMFGhQKQzUXI4NXEsb20l3vHlrJUffTpy6uKF919z1EE3thF0
EEZUm5vjR8iUsOjcvkPBnLVJKGp9s9rO1vSUo+jXFwWSbNNhyDO2ldGqwt6idBT8
bKgy6gWkzTuKg4fuKdy877Bzm/VRK7HSrrx5A/AwY3U5O6IeH/52r8/1iQzP5xKd
t4CJl5pWII+cbyLFl3CrHO4zFG3z1uxzN60YIw8P/mlVmZCwBu0RQh589r8f0XH7
TOQeGbFbww7CHmroqeUR5DzX/wT77Ax86d3SrSxoXRg4lIzNYHIUFFBP+yO/memz
SjWOc8qtIQEBmw0fvucQY9Ex1aHZYXIIdNWrzrZAKfWjEkv/Xz3MPuvkxC7huXuG
JDfy3k6jFYjxl2S+X0GqjHYGBahf+uBKyCxArfZPRyqPnD4TYg2sZoeey8hBUyPh
0uH3nuLz6sIqx5DyOm7d6I8zGlqL0+mOPqDmRiiHBF73M7hJVdnEs7pdeNM6aTvZ
Nz5ZJbsi7BHBiGT4AE3+zlx34HuFBqYNoCTzFEWxiLimS8DNlPmPOmn8PW9MHmXU
G13J+/yWRjI0b5EKpiZ45Xb43kjGr/lsLVfgAxPhBrvXAXqmqDRh/lv1XyanFvRZ
g+/BTv0ZBFGr7AaBoPa0N5ireXHrekMVjm11NC2TXgKbP4l2keHo7s9sZjl6ZM5B
hnJJpfV7HmJ/KTb03tUm/l8p+uw5CzLEm3584r/cEsGdU9MusnYGJVA+xGzhCG20
8MMT7FoFWOBBlkCAMV9AdG40WZwnfyr4vQP+/lce4D/xHjP3FkWWAB3xoYvKEwKi
bVHHlcJaNm/r/ZlEiHVog4VB99UQnupw4UyDrrEjA7FdMHmL+2oGFHEe66vOI9vp
b1EBgkzb2XH2f7bd12GGuMAfTgbgJSZ+YS2nysevXwwcKDlK4fXx8J56gqfuAAXb
ehOr7aNe9W7BDJ5Ut6LJvKduhPYU2bqASjAIYV1dnLW2e3mZ0r4XkTUGUUGfDdO6
8UTODFFCW9KF7Bqs9RKkq/f/lesKz3Jt8gBi0GVKqrPZK4LyWzg4DNlkSRmbvfyO
oBQqXcQVKzguzrK8VkdbsLvsZCdvCfUD+15/4y4rkOLu4dvKkIDdwKIeYGDNRc7l
pAyfbkAsqnGV6jK+uGn3zkNlPCCdsEVsfBfheuh7ZCdIvhPrKL5h197kG9Y2C0dd
+4sfUN7JK47Py5YM7gKXI7Lb+QawTblIqDjHEs4a8lSje9+YfX345jAjZW8lUD4h
JW9X5a+54Szp+j+eZpbYdrstvMxlQ46U+qE5ThoarRxU0vFxgi3UCP7wnrOjShM8
yTUhvGjelQMZ377Q/cA1jFMXedGHZGAugYOKXxBTx0nmE5pbmd7hNBCYAJOXt4TW
pkuAH003yGtk8MshKWmUMrVCn2+49brzlCrKZNniEkZ6hsdqeSk1SkfditwWBBOK
NiQOy0nSAEFunq1skHu63AwVOIUTs6iwqYITGjCNwnx/AHQoQ0CR73AT/OMRmEAi
LqzQFp9GHDn09r4wEVZERG/fjPOP088PjGtQghllJc1P8s8womgJlfPONdcM1Y05
aFIEZBGccuzHM47OyBbnAgxpY+/LB6jc8Ke0MaFh+89NdRb1/PPy8XUyNkNTjQZu
lsI5K5INE0yyQJTt2k1wgoorj8m7hqdqTBw3jdulhbUbuXG2IEiIWmrxe/eIZ7ej
rlu3Po55RIcHxXFFJQ9cYSr3Bx0TPPstUi+DVUkZ2huDDC6lmruhXhTBLWTLHdwY
NxvKnf9hu/plv5NThRxqZn8maFwJ1HD8esJdU1FJM61ByuVVxinKqvxtxPkTRPkQ
Cw/YodMdFSVAVNI7TPyiPT28pda0cWAXhvTJstqZk483j3OeGqnh2+dyb2URu1jx
Nrvhl02kcYt75+IhzeaCSYHrgZaefcnM3nRf35e8JScBAJOvXtZzXTICn1xZo87V
G2WcehGMwY/IwKdMq161VoUmkUiCw4c4zEKXEfv4C+lXtl2mCnMHoCregvIXzNHn
XyVAQmuh3zcoccq13a+cqVzZLw2qUnj2t1qcUQZTWYS4Ww6f5kZBTE/LUgbkbDxx
9T0TbiMZTYjKYaSJYij+IeJn7zwvrjNjdaAQ+g/4vBVKHB4Ms3BacLUexqNxvcbr
6nX9X8qFYD54yX9CMvfCtMxt9yCJbCfYugIvl7B8/QR8XW6a5RXWj3tb/tjg3e5O
4QTlvOllQl2nPGrExs8Qn2/bllrkXGeGrjERP3c9jN4MJ2IOveA+b4unSbiUS77t
OYVyi6MrXaGt7KGjIhklvBhjTFrYa+dVDvjYcT6Ice2A5AOEiDOiJ5STjjp02C0F
qprpPnOmPaWALnp1rL0R1QJ6YWkwD4IeS22/DTlXAjLRtX47LODR6dswsXPpZTkG
bfR5J9IpQTh0e9wF7KLFkq7xwq4bKSt/oF3xX5t4GLzykVKWsturOvbczGQ8eBbf
mPhknxsR6Zr8SKC0zkDSgCLb7d3Goi4KBpdR0daELkywcC9kwDEEyWPC7cr9SXct
m2cy5qQ/zRv6NUx0bZPdEFkk08qgtImYYlcoWyAobZHpIXOVKOQuevlrUMFUmO4N
i6nth2h8JZKFe3oEyzXItfirRFAFIDBdhQZA5EvpFt5a/OAMh2sKBudkAnIsVPOZ
qRvGR0VwsqNdIt05rh0HVTGfPMZKPAITdD9FM9OTDV9fYTg2RWaBWppiGuCfrlsK
VAd3bhxS0YmCl8jtGS5AtsmlWavxbas29bGlPpTkuJ6fptPvB39sXY0oaSCX0vPp
Zjg72pCFTHkcbeTSXV2DxtPmBZj/qUULzloKskZFiF11GXFrHwb1C0TacDJ0ZsYw
iGK0Rmm++EcIzcPPlm+sFxMpfbAVnmq8QvE4XqwZNajiw3cbjWb6UU85+zFMD8fG
MGCB7WyTKwFgpx8GHQN6dXa9xsZ50WgeGqKWRh6wzRtvZ5a+NWBcyDJkYEyNvKyB
bzllNVwz2JGR6jK1VCJKoNHTribjGYuc/VXLFARwf1w02S93wxddl+FdhinLtZ0A
zNI4IZrusFLqjjYf2iKnxon/ybNk28Wemp+q8W4XjUdnKAfH/UhOFptKDFdntcJs
qKnHoIe56I+nI+llPLUP8lBBTTlVBK06Q79LaQ8KEuCkXSTithdve0TnkT6VV92S
hLnUnESRC2XAAZ4Su7yrswJ2hFMVd66C0KPdTBNBTZrRe5xqEgo+F1EVL4I4vi+w
lv9ewHLBSh8m+q6MKR4Zb0aYMgoEDM8/hOG8rEqmJ3ukdaHTFvWkRKhJkqGg+tTW
zT0xkml/Gd0pMPl8CjT0LkNH08CX9I8dUS6PyhJwTrmUb/5BA72HSoqvoNS6/64G
hpVtceWRvnEmxq6C2v1Ems5QuN9JtGFL/2xW/M2iL7L7xOGlzH/4tqXHQPujhbK0
GTtf36K0HIbYZrufgogy2Eeap2VzV2D6jXJ8YIargVPrgTrJlfQ+jZc/OzMjxs3C
HbaJFEXrZG1+fDER29ZoGDowl+Fzko6e7vkIGBx0EAMAyLYYMcPvrcKI/JYI/h+K
d5vqHqjDmTEFVPGVK+xZENxYoHXozpIPBgCRF0qAsOWTwP9P5UGxd6IyYTyylcZ7
5MXesDyoADi0kcVOawgvUmRd+c83OndcjJQsMet931mhD9nt8ZlN9WrFuG61R2m9
GVQnMvLIDTvUCL0zBb2VW6sTEMfq9OqCCIhFSem0UG69y8Ow+UazZnzB6mvjTEx8
poZN5gEpTX0BFuzxhoqxja3oHif006PYsaLGRPMSF778Q7jSL8m4Ia2UJPSSJ2zO
+gJYa7O1lVg2mvkdBPMFwz7w5ubqHyAdIFQsBRPEDIL0Rs0z+fMaw45QHmY+NxWV
5rsjzwAeLeBG7lGlNO5bytbOWvuHYyU7C2F8EXQ4s8K89OoZzIZz+WDl6w7ZVDVK
jAzAyn67xpA/vV2h8PPxRuMGnwzq8H3uo7naIxMazIyNta4gPMeFu/O2jAS/Ncf8
vsWaaAxaGR7D7AaZZdbPxdF9pUB19/eizyFo6m5t3doTmyFQWui86H3gD6V9gu+q
GDXx8w4npMv3KEETwCJAWhIG3hiNVPvm6IgsWaPCeCYZ7FqCi2/opbhrX2BM6OzP
iB2x//S/7TCjle90Yq8qSBuu1p1KvsYzY9xN08brxUrZ240Rt7aXMGCaWbsz4UN9
sVYTDi/h2qizkGh4MwWAiuHT9kkcM7fwaAJ7QhQqGfQ1n5cMJrgF3oU+3W55noaB
caNBuzuN5Kis6eRUpUh5x5eFQs2ThAsJQ4d4SpNEKaVwLpNrVs9nc0r80KjGf+z4
YnAK2G2+08OrjBEUhsEUaD1UDJWmDrBXdPIhZa9fvdOuZkz7LjIRvIDRTDXl4ENY
xDIT7JEMNEc8XqFakgMwRyb1PKojiQAUxvfybiq2ZuyZ2Ew7zj+9EEcht63+mtO/
aWLOX+nwtBm1l93ORF7Bbb0jgJR0NidNP0F9TkjDv+MaHLRrfIzcEEJ2PoYlbTqU
uxGaGyUmMkfBVwx7b7uja9FLKL7TT1BXrhoGiwQCbVY+CaXsi4ZygqPqpmELIstU
+4A3vZsu4+3rzLZ2RykteHJ9tchnXGKY5kASqUA8kclTQ87WWdo6nlw9g7g+k83A
D06pBG0rwC4c5rt5Uyu/5N9LJBY4Vr0GmMLr4YEz0B2lIHkSXj73wKWAubj8CI8V
7xBr+ue/D3VWlYcwaLFNrFzUFnT45EWpddqyITtJXXJYoG+2Olr8AjN+05nYcVII
0YhN2fXUdjM55OEWw7e3Zk7Ws7JC2MMdyEGuwLfj3TFVkroi6YqJy2JbH76M9PyR
rwyFzQkutD0rQiEum+5eRkiZ/2O+2cV37AsEHZZgBVpwZZgL0HMHZXICtE6MCYgG
5G3mPI+T9ImV7vuhHOUTtjEnWG01yyVe/cmSlJ1+Ob1XfE8EZfLOFTuJxN/dL/yR
DVOff6sZYYPZ7UsZCNEUAAg5bzKqxEMKq9hEXcrA9Jxpw6C3gF+T+mAmmmFxhNtA
dwNX7n4ovtrhzE7+5Dz06nowS/tiJbDEnJqXxwGpo7TVOeBU0rNnfv+Rj8sfT7Rq
T9ilKsdFgdC3ycl7+y91VYjT5XVNS7I2wLI9Xu9Bu228MnCi/vHE6PK/4l2CwglC
SKxqGiRlJtI79sGChnY3XtB7v+8bsowWiUExO725Lc08zc/9XHTTYK8ShcAK/a3V
TsPoFm5lmeY34ZhMHyQMmVFmv4XFyv5BSPBD/eAo5pg4g8tfvEjT/Zd6/Cv9SUdk
pR85J69ktSKuh/SKkJxTP/coLieWG7TknuWNB4t+AmgahO1SUto2rbgkPeCs8NZi
/FGRyVegxjATmtnmkhXq+CtJVpFnrLnYxAmd0r10Vwro+qoQo7OPvY7yajJ3kp3b
Se0C0YKAUgPDfzC4FuGJPYN8L2SS5+WOBPcoeMKYErnk4Nd3o8iQzEgpvOWN/t+J
ngro5AoIpNy3IeF8EriVIQcAbCOJgDdcMQI9xHWcwZQq6e1Bdr7oLJqE+g2znbir
ZDNphjrKsVX0WTfTq7C2FzEG4A2gELaZdCZvuNF1sKFGdQGw584DnNEyleyUb1ZZ
FTDeDkADtWPZ2LknGPOzThfPY3z6mO74UkmOF2aAb6PTIRLCBENlADFduE/WiFwL
Juqxj2FvCcNKcgdchhIHfszmsA+6OZ4QEjdON4kG5T29iUKUO66KCCnLam6RajUt
TrsmAbOoc9g0tZSPfDJm4704keteKsbLPlQ6Le4gmtOxCNtp4kw6pMSGyItBdY28
TPlYhosJFMDDWsaR2ZbOKh90Z/VllOt/zrAD5CmOn1AF4b3uU0f6HGyeX/UZ3g+K
NePF165j7rk0anvLXYSoK4UllmZajtCOxGLSjtfP9zKip3dlS6kr4NUo1KCXUHUU
phuLKvbCHDRwiUwxUyYOCTyfecFEpQIl02Fycgze0zmTmYxgYB11R4rUMQl43Rso
dF488NJDa5haF6zG5aV9Xd2K2rNKG35B6p1/sidFylgE2ZsUDOgwakhvaRft3I/n
8alKGQQ3KxfMJKfTu2Tu9pXGxFVXKjox9LAZ2U2ZNBQ+v6XFeSknLxv370L07+Eh
51D1ZhyhUYM8oDjr+9biQ1BRIgfVQKPxdcBcWoYGFvqE49wKusz5s8LHiID8Tdci
VgP3Sb3tWy6MQjlhyjLeqTTbtMO+dKrhvL/Fokj5xuAHOMag9PEt8YbqsvzOKsk2
g6oOWDxsV5+jD+Ushot3zV6zhOMIPbJp6R084wz+dL4wNgPCexlbf5hohYRnWj8i
9zQIKPHPvJu8xpfaJSQK4tNK8Qt/v6Ua6vcu3l3NzxjraBvq4SSQlOLRgR4E4UYp
04xik1hywQFf5N09xEGPveiWOIr2Fhv6+Roz3+dSTL+B4RBKQCQKxeuGsuSpT2h3
LKcVIsgoRR3k6eTNLA/49+d0BgIXcz6BM+G65+j4KDHsfH8CG8m2NP8aI3R4Ffm8
acRruOJgXhQ2adWNT1SdrTSV0jLd/nBjFrwKhgGBBrUS5FZBAf9YaDWP5WYlvn7y
pqU0Wz+iex09FziQvQnfuY0Ed1K04W4mlzuAMZ+yKs4xOcXpDVITW31cOzZLi5eT
KUjIQTE8f6cfrfuKb+jDf9Dr54V6Ab4iH9nvDB7YZKbmfQQF+le5LZWYfjRSeHSH
D6LfQnnH16EGnv1vO4PUVim4cJkQ14BWsdrWdqEJPrwtP/JY3omf+Xlq8U4beeMI
6+SYjZg7OGJ1wANPmKC+Bh34c2edOor0l6T7lGRGEX7h3A4I8W7mKZI9OVJnbexa
N+44KcLKasrnXN/eKvhVv+dFC6deWqhjVMLJ2DXM3eeYoqQPL2hVJiWIbhajq2cs
RbaKZia7dPKj36K/XJKRiFkUKwf6v8XGJTuQCZ1dQoEob7T23M8SMXuPPoR14Lqz
ryuEC3uUTfHGQMEEByS5AS3blcZ2reKeGPYhx87KLdnk39/heIa6FFUIJX2Vxb8L
inOiFg/e+WXyvyADoScvu9z9rUuh7Xiiish2ENRsE3Pwh8lTjOgbR/GX//7NT5IT
xmncgoOCEzSKjFymeLsOjMs9Vr40vy5BV9CjMSTKMq9mxMurHboQ6skipnRDL0hf
Yd97O7O8ty861W22e6IhKjb08co+GTx6FIH5dM4sUNSFwSLp8WIDUGeyLAFHhb95
bnKfi3XPqc/gluuC/npoPan2Emfd0jU8BAK15IGQDWrfkvk0LXbYVjlAtA57Wqrh
u5D7RyJ4QHk3Yyh40hZ5ebPhzM1oAkgMTIae6LVGoL+LeyJ29sELjrNhTXN5HO7Q
LQTfuaLWTE6tnmqXYt0AMIs1r+h1MTLPvML9Rbe0NgeJWJ4N7u6DwoXRa79GEhTq
D61bnD+V3ndp6ILu9G2LV5z98GOUdTrIvI0yge44TN5/3feTcG7iPYhQpAFrZN/6
zELKe8Q7L90/25dVg/+ndp3D8EcYjGngevlbhy0JMcdkOdpsyGttQXu2JMPnu+6e
i2yTx8fOi+4HUOl8CCeOnYJWSvTfPcIHA3muIaRawdlxpK3Kyv37x65A2tz7rMEt
iTaQQRqpLmkrmlAdZv1edxrgd2q3RoviFy71ePMJ02x1/H7SMRGZCLcwfHyugxuM
FpqxWhMa40ZjUlG4GyZqegEcVRkLBAAXFHRT8qLbnyvPnaShaP0rxwWyPkQ7ZqUL
ebth5cEwa71moev1za6mMzRg7CLD4jriB60GgWphPrziVWSmgPDjxLDkZh2dXwa9
yh30K41N2bohdbe6IE8bmz2UzuXepK6U9xQdsMe/ytxF/elhNvKP9SRaQe+vJKDM
YRGGowpaDsLEUOcyHSasBE6m7KymH63VDGTk1dCl22F7ZEgB3nPw++VKGLhNxwfq
4HFEtx+GiuFuEc7mv6Ud9Ve6J9VPWICCc32OrAEM75GGRzrCub6aZA8S+5tBICfl
ReVLzPjUa7QhigNwpLQthDpsjeNOOQX0wUK22uw3kzPtY8xEv+8RZ309ord5Jz6V
zd5glV0BRR7j9ys/hyjHNf5xAADSNy4SYRQj6r36t2mePoiFIvG7Yo+r5yAHsyZl
lIz+jzeo4xATK4WDNQiUecQaHeRktvv1lCwevfJEE727mYv7PhqtlPtlKNHD5loE
lciyeuknTD6E95nON6O4baPF432IRyEevDxhXjylHchxYrwfrNNB1hbYwhc/9eis
KOsypeMOP0WNX/15zyirND9McuLIDbck2PfhOFQuN547w2slIF5E3byBlaUZgkFc
cEckKUpuBg8yJOqyPAET1TxwZofbA6Z+NuAa73bJFX/5u3gyH7ij6tr1QuplceZt
A03v0AAx9Ss6LonQKCXVdq+yg3Girni17RK6Iy+UAdIgvP9qmyFgbRneYsy6EgWw
uSyve47laCeGYHbn+fuUWDCuxlHRIixoSak9OsU21k3AdmDbmlAwARS0AVPQq95T
sKc23SIgozk1al9O8MNrNM2AycMe1z7BERuAD2rBJ8e8z2eyT2VzgkLZB97qKABL
37XOgtL1VwNMvi4/YRjceADz3VfDu5IEEsSax6DVpArMgqNFbSxVycHR+nAFTaV7
wOYSdB5pU7eL8L7sKNzgkDt9fKNAPFFLCOa6v0CfpdcWjwzhX4bxvzlSBJIqOr8Q
S9UOKcNti9xEgb20aLC81tJpZTMGpMp2gGLNCkPXsK7AKmkMZ3Fji1tfYNp6oMkt
Kqo2yqVP2MklfBQDmWt53AcaOrXRfq2sJqKhy2wpFzU5oL21PfG6W08bX+ExOX0s
0r9gJVJm55Lq7zzMC/xuOH3FwsFafZ1zu9FF4rMBJET9UfaZkSnKkQtkcPxgBCye
fLQKGXXYLhtdM8c8d6kU0SmqlHoSqwBMVpaMnYn3CAMEcMpjHYa/6Kcq1w3mstAB
OLlChykP9NP3qc83wOv0AjafCE4NGpuT6x/EAnAPMKBhKkLTRbWZsmDPv1DnCd5j
GNG/elkaB6UfpNdOqehFoOt/wywo2NmFl5q1Jq6YE49yMToFphPLi7oOw1oSWJBF
Pq1qQeBoD1j9yE7WUU75vybpatpkaanf8xHRlmpqDP0IVRXab8PcyTzD3QTkSXlr
+1jOz7nSVLtupFja/OefmRpZKTPaUNhvjsgX3FQKOx1x8T0LFeCaq54qMvEdxrT/
bue6m4vepoD8ayXH5CfxpJu3FxehYN1ondfIELvRCc1FbMMNfRIq6Zk+LyVO0ftz
kuoQVfQyTf8oD+rsn4OURoWAW2Q/h+OMGJ7fvMW5UOZn21TkQluA2I+w9OC04q1E
8mfPZyD9cNpGV9eCzIU3MNN1WlVK6xiw1z7xLY40pVbLQE9/JA1d8eaWWrVSMRtT
qVf7IDt05dYC2CRr3o3wynVrQrogJt47HpaQ67VxlJ9tHMGwtiilcZjG1Djz7HDY
2eMLR4cdKVd49gy9dBCa5Qoalzy3Wo2DJB0tN2Wo5+WiU5ERSNCTWVwnYkqOaatq
iAovIMKg5Df1yLzwPgySKTsTvkrCfoGj4xfHQrakPnYPb2Pzjq5rpoJXL63kKgQn
mJE7R6fVYTMpIYY2TXzEy2poVD2QEAkEcVIu9WTCGP5LbTeHpUnXYQ1h8YvpRxWu
Lx2NruxFR7QzUIVATcPTGWGXRni07LbRASlVyc/QQfUblZfu2hKj958AlSAj7H0p
pr+WFod+dy8A5cCorNPhwA+YznAZ8MdHTdgmwHc1HGMRlb0khUFU4wdbQiAqRIC6
JuyxM5Cea8wd018PKWq5W1ob5WaZyTwrIdKpwuPxOvz2LgTNpykNRKyew6gKjCvZ
oSgr5LiUST5DcjojH5Nje9W/Urfgkf+6hB55EN6KW53v03n3rvNuBSyf+s7Rffla
fmSXyQpZYEiimLVQAb92CPu67AoLSnXf6csISIqQ4osmO+/mYyIy5olFP3vD5Dpr
NGHXKlMHldR9AjrLZbVjXWl9V7qh6FmRq8fdZ0TU+Z6X6U1MUOUVlDtSXEm6qY8F
/ksHvwHhAKSCKKW/LP0a9mL6YgAqBrEr+o1JaEPGUMDoR1Q9kP62SQoxkEuMev9i
oewaT8xuedgnMgSHdsUmLeBHO2Z0OyzXZQnh4LB9bDyEGi2plIwwDm/YOEKld6tg
TTbdjNw/GuiWPTx4Z60a6zr9NyPPaXPKOL5NGE3vfb7TINfrU9G2Bd652Ojtdunz
WwjNIhdxvSsCcHKuAIZgSbXrSg4K2YBeCxL+SvNhWMD8WvxTnpaIr+fxRqL1lgjq
sPFLAFtqVspMmvCND7TaIEy6FssPZph5etzP1teN08Kbh51AnfTgwQ+Y9xt9lGhJ
lynLUXlGr0RuAGSD4H5FUkNyrKLzdKDtDeT2PVd34FivsUW9UTsFdeUQSlcloArW
KFca4EWmOJT0gzfliRr2gx8wmktqwW3Ez6zuDbEsQ9r5I6Y20BLi9c5eQd4+mADY
Jt5UV6z+E8yj2W5GLVVVq3omFVWRWk29KWBfu37G5hpWKrthOTwhwpQxkSVNR/rI
/rLWWbgJyB2+jwjIDMNsk0XujYBYnFIFPEqay2yDWS8p8uv3VuHBobS0Cz+ajWE/
2NXmwv7W3IMurvEwaSCF0XIuXjKZUu7Gp7TuTChNJzAlZRB/hekPjEwzMQE47Ey0
vIIEGmjL5rxciHr2lUi85I8tXG1hYoM9reQw//V19/lIK+LhMYgMAono5IZCz9/c
yV/wE8Fi6l3NxsIVuLTY9GMvnN8GgImecFspsTe3fq1HiIQNZeVw+UPNjfHSQDYV
VaLgPijqQ3Np+BeMNdCB6E3m6/AcXNCxOE82rFV2sJpbXsVPBXkhZi0U+zZ+YO8d
VJIlMicWBcpB7uEhWdRknuHNTcfSwxZQlsPu7QekEMnt3jv5s0o+l6XA+jUVb2SE
p7jLNS6T9yPpH4KPsQRIhfklZ5qQGlB9sheTXmEUP7sxZdfP+YYjK/i0O2XhBJQv
BQOFwrHlrrRBQNr16hgfn3aeHsVeLKY1+8HgzVEVrbFYI9+R5VWsDiJj/V5XemCm
5ZSXiP3K02x80KqUNAjhsl4tSoEFt+F1B3OvPnYPQc7qYi6ksGZk7CQniFAC5dAS
spFZTPznq1IXe78kzaekft7BgWKQLhucEzRLhp6z4wKMX47rTroFeNrwNIZdHZTN
GIXmkdr8H+f4D5bmqBj7fhmnwRYTDiAnM4Re7Nup5FPultJ4GtVWZxvb5K2Cr/Eq
nozddl0L0+orsArTlw/yWLIzKuEKK9rA3Tcq+uG+0GxDLyiK1BjdJ1MV/OGEAxz9
6CMMvzArygMYoWZ7eXmUCQz9jvlJqjkXx+jBWKPV2Bol3hKMwATrUaYGdroxNekz
Z8BusccVaDZkxZ7nWp4Tlg9fsle7Ry/Ium08nY8+x8jrNmE4pa/nhh5pzK+6aMMf
kfK33Xbt8627S/mDoro9G1Y3Y2DA1+PViedZ8sLpoIDgeLAxzfY6vTfOW/aGsJmF
CTHBSeSHFOtaq5rx9mKlO25/kPaqBhgA6vtGYuX+kpDRd2MiDTl5pG4KM39gve3k
pl+Zh8zIA6DOIasL1pnC8oE0Vw4Nd781kJ6QDf8EGTkucvYPVohZtDsjWv4gtf9i
g1rjrXj3StMo/9olo/NNCzFGXbIyIX8W4qsTY3noxOhy+MbPtUV3WgHLk5Oc73dd
VoA6+MMZskuNUIl0GfGSBUqkFVkpBIr2rWGoUMtnk5TV2ngAdIQpJ9p4UlihitXP
muDZtPAHIjASCEqGf1+9BfAKsaOpknppuRdMm8kOzD0hCgauiGsBowfSSUXm0doB
5NQ2k3hIgVnUOGRDwt4QW7e0dw+NRsXfx4FOzpiCne7nSBE8eVRrZ9LU/nv7yJZd
1yusbeVwEw/2KVPpet8scUCo6kgV+b70oDO4sOqslBF4iGxFY3QH/mhM2YNOwhvu
X6EsVVw5f6MGPAPPw0MAHcqQ+8WDeQKh3rWNC/gErmuToHKwHBAfqhVPQI7HXWPC
+Z+BR/MFR8VgaBKnnstvNFEkzsD5fsELfdE/V2f+H+OHGyNNghq0x+o5meAhz0us
RjOsxRKs8DK7m6vvMPui3y8v5TO3Wp1YTXeYiROWOF95Nzqoyl5nM1ZJ7JLDJfrm
BWA5RxGapC2NE/mdF1rFbbX1nNgSIQAnVMnEpkxmABw00VeZfywS65P5q6BRpONt
NO1GGfby6+1f8eagbITmISDvYyCrjH3Uq2nUooFtgqT4oUgrsstXCCCa0/hbSbx3
hFn66AwscktPKceU6uAKuX2oMqGZ3jYjW08pRkQXoVj+snzEO8IWXu2o50ey6o14
i+b71Ufc2wC2uih6bzQMdnLDbjtdLLGJiGvPZDd9lgQifOAcJyXmLsoEWYRqTH9h
Mbk1AG2ap3N6+UWYVVo0QYOoMZHOvU6kPU5YkBPLAXq3WUAWrd7l4uuUvS0TN8va
JYB36ecsiHrA9nARZpFcpn2zpIExbHK30eTjv8kP5mhwxvRtY2x0pYfcx6LZsFkD
zEd+GU9mMtIAMmhL1hmDtY7bJKSy87+EOtwHJMpFrWQXd8ENyb0CTQYBcjcRRJkq
vKZCHkHUnt3A+cdZttj3JJ3mZQBoE04h1uzmL1UQbxe7EiuCU9xbiHALPxoUuHNG
OcR7+onL+L8ZpUDA8LcKdmAgm+6E/4G9RIip/OI0EGzJt3WiBJD6sMEXHhKiBHpn
Ce+dvhs4RcPHrwr4CNXcaN6vV29sGDx8jNcdLTZW/4j8AEDQyLABxPcIoEiim/TK
qdiD494LobT7mZO1coKpsKbe6oUUaXd4MGtiyUm4trdlM+dWe7K12bxj22yHpk2w
nomCQLraTF0TycmV2E/tOFaGtzeD58gp1IU+oL5OHxYPBcC05Ksba3saMK7aRGbT
bu6qde/qUlGKekWmFKiORDkfcrhInPP6RWvsUW544GxLYPOgkX5VFJONbV2NbcWJ
5Kr9+ZWwx9kxXpQhr503T2k5I9ytYD1mtpTRswphHq7zPfAl8lpSOX+aQA9CJ62E
olhx81zgSAj5voPj3XZcSA3gDv7VQV1bVhpbenerAaMK2WeuqbQaQtDsI8tmfP+n
+uzSA1+SzSkhBvX9GyAqDVGErXy9QnT8IUNzGZWU3gjXXr/zo+a4d1GtZ1gd1Bq7
+KjvrnzY4mPnCAoiEKCymRBxbS9DJLMa6eZDOrnLEB826KSet0jkTKjCbijt5/ZJ
kLnM2+wVl8UIF6jFumGn48VpSFuhXZWSUhCFi+ZFAcNXG8rw2bRaQepEkcNpSLbM
W/yTYrUHDBS6H5wNhPz8I37SJ5tvOlLXi/+9+pi9YFGtansBke/RzD5fyxxEKsJn
xxkj7+aE3Y9NFGZp9lyzTaCp4e9DBXydyrQDqJlB+kGVtysmMcFneEufPczkWC5Y
mrJ0aObug796BTqeobJoRarUeTv8OWINFGscYj6ZOVhqgtbgRRVimGYeGJp/OOkN
oF/3OKY6CQnTcGCPXbn+QaLzfnqb2d9mvHm11/5DiLEyFk8bNkdK9b9rlR707YwY
mSMxDzxEbEmlTddCdlFMP7bavsHXEqNPBMH3eZdBaExCuox91f+LWYhhE5m8a6fR
/9Ec8qn0K1VEZMxRM0sK7wiN7N07kmvu4g7blVfre4UPboJWMoTGZpyEOIjSMd61
yJpjB0f72ql8dmriPz84okSMbNWFdAuW8ZI5CDtO5nFJdaO10eYePIw4Xy7ugKsv
vg7HGM6A8L51U6eXOw8OhPW+LSsAElVGyJ4pDNexSDNw2wSEdbwDjfnmGs4KrJuc
Na0UeDhDFwaujLIfb6ENMxxUP5tb7ca7gbE7ucjbKEutHO8BfNqAqkXF1NL+LYzf
s0236C0kb1QgNsvBQvF4B++8u7u/ul7Kfe35pEIws/RkrCVaxrDn7jL2N1sUuO1I
g686kT84rptdOLTrTe+7S/8hVaMdY6BAqIqbSOIqKFOjzrJVm/VCgggQA6OLzckg
ilZ91dMOm+aIuRE2mETTEttkrEZ6W2KLV2m9SJyCxvxmy7FHI7wwWKQnpZGNety3
cWYlHHozYUMBbHJ065/AUMhpj8mSRWwsT5Wd6NAVvpidKWfJhX+o5dAtKwm8A7rc
KOyPK8H8Agsg0Zuno4UH56oN1Wf4OYOw+LNhutyhbQrmhbXRl7cL3FT3nztWQqiU
Dtqq5BOVpSlyggCNO9Th7ihDktUMBwktJoVZdLwF75pkFfYqTfbZ+ak62aeWI137
sbXc/vE5F8g7czFAtIDLfmzAq62Xt8mZbIfHFQxOl3681lQvgDBhn1ua2zBmZHaL
1hVHhiur3EmJu/3LqiOyp3YXUqgCErSztO/Y/4d0oecbv6U5Z4pz/4H9ocZrLv8j
WmhSSZO/9CRJRzU/2xvm+FvVTW+4HtWHNZcuKWqOzHiw8ztF89lmKqL+RFWshFQm
CU1PAnTU7/dxNdXe8NzUIDk5XAJoSNkIWxgglPkLDZObcl4V8n53EIy6C/oLTrg+
rsGNmbUM+H0RZbSQ5mj5sRMGSYj0buenP6O4hw36xDa6EiF705dMEWhcwdec6Pgs
RZVbqc0VKUwTKvainBNFmmRV9tGIQ799ZnxyZC6g28yg10o0QdWF3kH/Jxd1Vt8+
U9RZc+mesvA389YSUs5YoBr80IHXWVYv8jINcdpzIJeQfJ9l7Bg3AMtQUzYAwoan
vTsrWWe/SoifCrTiS+lA7m9vrKXL/cAnKFGAGjq+JEyxkjxcxeTeQ3xFACgGlkAl
eHanHCv9hPWDE3DR1IPRmceNC1BIESA6fRsethmaTIGZbkWMHTjOy4PO4q+O4mRh
JYWIxzqxkTgXRDKGuk4Cmqd4xm2gbUB+a23TJ4+1pAQTcQYehWZMjBS3m2rvz0wQ
FzjvHpDteExdOGeRejI++3MLW3jVQ/uucap1JywSm88hZipb6x8pnzbHGncud7Ux
tPbflRzZ9uI5ek7Q7GUJI9NcjmPy3HKYCxJ03DPIAiZSDs0zRSdgGlXhL6/eLC8f
UN+bAatuFaEJhvyyhVo00bJ/LzRi8dMcvlk3fiGa7Sj95JOi2KM+liJIoQI0DJdy
5JCEo5EglMyFrzaTxcZBwWCLvoY545ISmgLXYa7DBWdcRuvf2Z9vQ5vGtpihMfXo
heVXzD7urwkzdwoz8a3LsyHdQwG7FjqjgbQor9wd5mfo9a42XOX2y69TmdK83NEd
w+biopF1kH0Tn49PUQCCuJMcsYDeyskrfqv9FLxI2R07qt2PPWiX7kV6K4+lOh2u
fGqCFsFc63TPEUc2CcEoZXFcoftFK0Nktr+s7+SPlGWvSiW5KyrChILhpSbjTFKE
uVxN/PbY3uvF7nxzwvuIn+LTWWpjWrk5FSMYZqT5kF0jWfWkG+MWEz3AkX1GxHUy
u7nt7eRcO57TG8oZ4aF4/eoWDD6xqzivF+29zPaujEmfr8vWLW7gl44S7EEJJkSU
1lKXKdppBLJY0fm9bdgSLg+gHegDBJxiOBFNeygcXxYX6JigyNWoQ+CkzJGBsPYc
ZItnaRyNBQHJb7IasgNlPmsJL9qyPxChaSzPW4jR/7L4Ny2bsu555BXxseHF5AcE
dSk7rPEjTopHsNJFW56gEbbnvbggIqJuBCxFmG+OKFqTmk4JGnI1Y8Yy9HWOfMpz
+WEqnqBT1o/AwYw2sm1FJjbKP8pc6Bi07DXfITFIKP6Bvt1YEdvafl08B3HeUq8K
8xi1LGv+JJSr0nUD4nIA4Cshl7nPnNlXaUhv+JFs8t6X6r78+AGLX5OHUT95ZBZ5
jY9XAhsnYCQhlGiZt9ScihUDeKZlMH45a5oxU87Vqn1ggOX+mdBxMbqHoxIZoufe
eFWdUq/2Kglx+Olw3cHyeqrAfVbMBbogrYdDxLur8iOccHrUyb0NyUngScCEltS0
qx8caoBS4X4VQjQqkAcnUFqdF1NT15vvVB5wBPlRHx38pOaKhG2GrvhUc5OQb+Zs
2b9gN/+ncCc/vJ1bOlNGUsJr6lCiIg7c8pZbraXYT0BT0nxZ4wNMbPhEYRvUhm+L
8c8nr6WGbIHF5MqZNIKbvqa1GvhV+SYBE0YR9qGmyU1szyK+kwlAtjbYr3ezYg0N
9NC0fpacgY4+0b9L+K5TV8m2yeXBwolV00HGlcQXQHx7rL68rj+FYRILkq/oTLbM
4DfvWFRlicfgWcqCt9R8sN2cRgi2Gu5MaBQgxRMvU66eB6Adglcsk4JzFV8kqa9T
op1OIgZh06O3UlaQeuXHvr2WyhTfFWmrHkVmPmUnPNxP8RSXHVajGkEfcI7lnScb
j2Kx/OQw3W+kOnY7DIQ2mx/kMd79IkxC/XTWakNKlcVX1Cgguqfb2Q2OpdCNF8yw
lEDXdutdy3IWqiAIzVMjQvmfyrc6CMg0GTIcIWnksyrErUseWIbrhHEgqlMnANRX
aqNQskTj4yxYkYRK315y9V7jQRphyVTR/ibVwQzDxYaKiKjC62oHR1z+lHeZJ/Io
f++U+/Xamcq5YVzcvkPPR2ZOQshjPr9QCtLyjFDJLfUwuPgYi/F8j0aBE4DNA2Py
6RqWE0wBZ9ZzHtIhHhwUOmn5aQquwsSlEvuFCv3kno1Jn+rakLwTRrQ79vjSb0g0
SNhyOdNN6ZWgY8kNQfZZDv+s1MVMEw44H3NR01SiDe6l2VPIOx84l51L7wlX17Tv
SRHJP7MtE8bzuBLfoOdVlFr7CFGrc6nuVZUV/jEUAgzOW+Z1urFJEf6MCIEawL6L
eBDLdQFydsEviyz/BeQMjiccasZVppQmmOP2cWkBISagtfUZMjycK7BnZBkamMKj
OdnmZN+UkaekUzULw+qGi8ibm1wiafwn+upIdLwSsSDstYidf6SDkPfZJRlEKeNP
EpVQPk1w8twBDGk3ReOY2ZrwbEYBRUXwT59IHM/CB15krm6zo1tJNQiW+kJfDnYd
5Tb4oKo03y4LTvucWjYJ83i5jmPmVzI7sFyVjHmEpmyuRnGJDRRHUjsDWMcgeNKl
oxMpLyuCF33rJU5y9qS4ocHaoUFX2HFYBjF8DpH4JN06IoEwOJIUrvVYzuNLjw81
5yDxITAxYbhzYRQpkQNRfBPoANuAFLztIHtyuabkOAsH07cBnzAcZ5QAex1WBil7
Sz4cGuNJngE7g32NhHdMBVZ4e9mxIrcbvXYl6dxTHF20FR4TVAHzFeDdsUup3tcl
Caun22ZnZvlaM1rZTGWRaUoVUFjheIm61YYCnwIRiAPxwRJ/ouGR/4tRLvRCGfNt
9e1OtyTjuhk/64kg8RWnJBp1kb7eJz9ZByHEoaYhnWwkksASwEtl/7bKz9NDaHFa
r9E7q7oOJAIMpCJiZiFVgIO6nubZI+b8Az1kOe52484httvGJpchxoj1vrialF5L
mrQ7crqmQCHFOesXrJWv2Ef0ySaFQF3cHF2+QIB7h0oolUIaH7/FL/FLqIiVNYrA
RI4PHRfWLzXhdcicAATR6QasZRnSKn96PZym5smA4t3yFMIk1ErJj0uNQD5KV559
bxck0ow8OpzuaP95EgmZwKufKh7XuXscEwizPn9mkLs88bX+JzenLusAM+9H8Wmg
DeY/5GgW/Xy6bo8nSbXEANJhx85PT3Enqd7K33ALyva8cOXiDjdGEjOqjLfuPpGP
BhYW2TCYPDkymGnOsszRfj9Zx4ZlEmRHuaP0RoBXo49kSecFMQYKdxTuvUaJhm1Q
GnKKFRGmqlp1SwYqk881lvRJJtSpNgHDFaL8LQFrieupGt2LSzm6SLPfG+o3/BsL
f3bm0Ih94QhnhxpHpbC7yQ4BslISL2abl+jCWsAm+RKsrJ5Ka4XL8ADYke+1mJt9
1DOa/2nByyU9My+d4F/d82+H7BpoCF16o8vjsIZG5flFxQMbjo7IBO6OHM0D2R3t
2/F3URLEwdSQwPwVCmKIlbgp3Ma61Cq0ZWhrnjWMqgONUt7SoMviwpHxKIYWGiLB
U6l2oC7ExvrFNePXn2DrfqaoNJLN0oKI/1MAW2mN9Z+Wp87NqUlUmFSV0EKSPtwX
eTUD3rz/WVDuHChE6xUY8sFxpdAdbsufATaDmrL07HBRL4OgzYOubabrRqVKpSR1
RMpWeK9GDgnlm3jR8MUvAmVhrVi7SdMKRVk7MIb2rmWoKNSwLiFvxKaLM7/pLnrX
fc0JhRm+IushuTU+tBf2SUmrSDN+STNS2QnJcbkvcw6XEk7jq6LEOAg8IfuyhS4V
BkXfTCYQhvdp0aV06VqoFWafQ8oezm/U2QbddDZ8SD1MZ50xuqOCeMBcQ1Cawm2Q
h5PF7J3uT6b5wwaxvM/kTI3j+PlGi0Mx8ycVUISzdph4l2yG/x36uxt0Z8aGz9eL
DcUUM3Z2Jl/iHPWhXqKOw06fSgEmhCX8xaeUvrRMBYZDFgzjl7XSezK7Bc0KRZGm
3MztHlm/V/hnp3Jyxtvz8bCX8Tli71mO2pw2nwu1rIIPDMOSzWnS1hXlJ4L5SSyU
p92Z1UnWMo6bvfOZBBxJjIRkV9+WbDkwvnES05ZrSv+h7iioqU7Y3U7GmJ8ce+w7
NKA9L06auaJRKhhizp9ZaZGg0JRRC3mk7I375W9aNN5IiAHWnhycpRBWtYv4eG8A
NooK3Lx0kbewXlnO99Su7olycoLrrRxTpvXp8MXwvbYc/G38E08nd8YMwiERaIYB
ejn1635N9zWhnrMf0sY9jG1a5eFrhDCwHPRDyJMnFEuaH7rg0SShXQWRpiEkZOby
miLsOirGX59Q0Q2GGZ/+o0lv78B/vfyqhPvPeSKAepyXL4hliFPrXjmXo760MMGA
eSg6zcz+xnn9ciIkmpMd+vvTYckKozRzPcYrV22GzhjEyr+Zv7qyjWr19/7/y3Xv
+VH/0rPKdHR/3QF1UxSTKCOigfa0UKRCALqW6PDhN3KDwPByyjNMMa2e2AnXc6WR
w5LN4OxmGLT33JbH5X7lKoCrQVMgiX+xyifu8AOLf6H7kY24DBLEMB32othK+0TC
r1QQ5GUY53nrtz2/QWma6AfdzSCJnzMxd1uA17PBz8cof1B1mtsRzDn6ILi5J6yR
dHymKTHZEXz8KDqtHLO4lykkCO5OKB+DhbXBpGx3OByRbhTw2uUvkUadoPyD6mG2
8zMusnPowPNRLm7oXvEEZjwZtU13EPo6I8IXfAIVY4ynTeyQsz0Gp0iSxGdu30pg
ZEYm4FHhXfHAQH/qbnuqPjhEBU7QTZRk2NNWVjjSDofF5rmF0RMO6Avq/9P1gnQ3
OG9YPRK3LZ0cEaFLafGr2dPB0cn5/SGs3Bokn9Hso1uF6bTJinRz9bnA6YhFzOGy
9XiWiNLA8t1A2QxkoM0gdNRQ2UETE0k9B9X4ohdHapBWRz+I6Rl09mMmKWLtk7HG
OLd9Wm4tPzuxF2Xb7uCcZnokJPXEMZZeDkle122RFMxvRXoje1LoW+724z1S0k8z
886kJMvIBXC5NJTNZPa905/CMYX55doDwjJg6GXwG+1G+tbAZYWnFm/125cpUsoz
H+T7pTnYwBG0KqzbV0xeBTMavyRDtq/Bau5PXHlQ8igPWy4OPvvJtXES05TxUjun
e5wWx6/myn2zocsSUAC/al79JQgRZPHDQOk+wXKC9M+en9dvK6NU1XlciVfwZuOZ
VTHVHsSUtWKbc6Ar0cRv2A1vNLWEfmZHmwtaSTsWPyH6rR4sQYPBI4sdpL0kpe07
nYOpNQzU323vhpUjUTWajpD9bt6Z715nCD1U0NoUL4nDKby9egCGrT/bZwRiltjq
slDMCbtDdaSIEa40aWrItW1i49cs9T35L7IaweNhQPZt7bg67navkXr8C5yC1bkU
cGFv/wSDfKdpJVaHiy7nXenHPD7Ys9L7J83MJHwGDMOBQ0lAMdj8EDxuY5pmHXpb
xERaP5TzEdqpsY3OonZKzHfXJR5koVuG7qA7DMjkncZCDzjfebiT2smVuac9l9Mt
/+sTcF3ZzILx2Trt7xXz5fQ+eRzUQrzwgXjEk9e8O/iR5CRj3r5D3mboujo+jw5i
DwTgoesHFHjDU4X+AJu3MdY3Ek8VRW/qkO+7Z/WLNgzo/jApz5PpHbf7M6y/azmt
KFYMfEqeJv28jGE5W1jREIXdXsY5Dsq53VUffOuukg1hhV4vkqCWbe45Dg1Qx+4T
fE9E+RVruTzbFBsRItWk30TZxYX/AG2dcKHyvgkkzMdMzw28QzV69UemkknW00vI
o8TQYmuLdBVr5n/cSN7n/izBfuRwJqN4ZzA+u450fZHoyytv76vgeq6/apMt5UXE
wURSkq4aNGOJ0JsnTUvIPyjoApcZNcZhEeXFuJiwHYDnumcYpC8wg2eYMGigbBVN
3m9okzvMKlToVUg7pcmPjApiqqGKTMwl9z1MD/oSTc7U9fVPA/P7ftsw+vdjF50H
QPwgjPSWbIrc7NS98bS+e3D9oFHCpKWt49L36RvkGwfjNdyGa6C5L01br0MT3p7m
2vx4N+Ke2wrVwll8fEHNZhkAjOdjUqxUPInHcuoZH1cbPL64GKTIHTwsc9UAmR4r
1HDKTqQDhXfVSZn1eFvsav9i5Z6AkmaosgCtS9+UY6uRLwStgeo7mcMZewVZGWAS
2hSHKw/zqf99anyEMdfcIHuObaJmwTuJ27bS2EByA9NWX2pDzlKesOrNZOb9lpa+
69FWTohyCque9kSf1WAdIvA0nC9XzC26oQzaDgulq7hFlXiZ9hlsG+2BROQMS+oZ
3cl7FYgQMIgRYHxtHzPw36aDFJTNmqhZekrh1ti8Gcyeerj/v7qw4XRxTLg2fSuI
QuSY0vVo2Kw4i1BzxcguZuLJFq2kSCAe8CQbr8rdqaJ9rBThjA6NT9H4j41gJAhb
iWH6ZktBBixGAUYx8UoLU9keIuGAfDKycQ0t5yyfXy05kF1PGVuPXGkXpG2vIyrm
d5/yAd6BYu9JT8hU+CUJjlu0mzbnywSWvlI+pM3ds3p926IBIrVwXkJdXDfuBdII
LW2sNjcDIxTf8a0GY6Hkx7+4GHVIP4VRW6Nibg2t1kFt/YNou6sXQFvDjz96Hhdm
hFE/Qsn3FMExFLAgUL3ZNynMy4YZsZZTaFqPIp5JKYZcYpn1Lz86kqQDsqo4KBlp
JMuTN2Fob/ljyg5kYS0fNEh/Itp45r1DyPL0GMGpcN37x4gAD5xPPi69sKlZ6sUZ
6MZHn1/KUlV6Hd50CQAnBhUU9sOVSSAF68ZHHXl2ssE5xFc/vgOp2N6CSa5jkD0q
qFHI4SEh8gQNgwIhW73eQlydn5DqDElm86Bl2dN/tdsrwlJBNI5ls/Qzfe52YIF3
ILpd5D6qC4jls37ZxN7Q0aaXhivRRcMpofoScYUlNP3ktuK1xMg5Nf/PUIywGweQ
ILN6HQtyWOe+p7lnhzHHf7sVQ/LB6MnEyTZ5PHPiLqe4Uq0fiK9hIV8th5wrA9Ks
3k+g0f73LjvxZHa2cNQGZ1Otpdrtwk//Um6IA9BLkXd+9K9gNtdp/wGuPjXfazsu
HgA2bwustnCMReKlRMrqEIUFw/lHEZneYlbVD84mncmdMW0ObVEhhOXj81sVi5HE
fZbkWE3CraLW1U2FHwSkAYr6HEuohZmWS5JGqY0L9B106tU4rjx/cof/9rYbzbGa
mBPEMk/SrtB3o0pr6fvpxX2AZrP6Wu5PQ6hvkWS9SNcpsQAfR1zhX6a+hIpIojFO
TbXnF1qJDXpgUSksOlKhz2FVeNJRY6HTgoV4ILkR0UvqlT0u6U68bynHEBEwK299
jeUi0wCRyeTaVVcHLN17NsUJokmUgi3GP2AcUbhaIQYvzFlIkewvuKxE44cSKbGn
J+irviEA6RUEzjnLTG1zyautx9dfBqJM2bRg5Yvy9Bzaa+0CIPjh5prD1i6TA4QY
zFRc4FEG2KlQFc+DpbeS7k/ZCwWdkBoRdghuPUytYEewV9we1viCUzp78jhmYiB+
N7kZJuTx/E0s4b9F7nKZwDBopLblcnl2WMFZquWA6oSnPnKSPLBmrwjirXQw+Gu0
TW7W0oxvh+DjhvdgWq7qcWhY/h6A1n+U9x8CmzrOjqaEhw7z8KppkO1TFEgPiWOu
OaimLkYZU2fEbQ6OBe8YQKO+DN3DpdzJDwLo67Fzq8ZbWAshzmfM1tRaDdqGqm4y
Zbo4HqHfAZtmcH1wcywJx12xVbp/90s546EbwIckwYqn3YWs0j6t1d7DbJHbuzsB
BSu1xW7degCHGG0qUz6RTamrdY4ek9CeyTMZyCKkh7NunWDwtY6NKFp3dxNdM5Wa
lKpydYgzFBuufgRGW/ZmnvpWrJ7cEfEApza87XzaHao7KqnH9E90UiLow6WX45ZE
iu/ACMJFKsI0EYZi+uIg6fICNP+MSr5IpJm0+1tAbUtk05z/zXcYSndv4TIRUTfH
pJyNBSYAumRQBoKGpDyt+6fFhCXSPsEQ5Dlve6pgHL3vIzjo5G9Z8cqujiOcPqkU
orAN240WichBEgVsloXVWGc9w+eXwIrUChNdTyM2CG/ptxU+qG4eiBfyZzGDMFtT
htJ9a0YE02SdI80PdXoVdrRcVYoPq7GnM0P5DABaGXlmJ21TvR72bh2oHzs/yhlQ
+XFYpKue7RXjQv/FL5Hwnf47BgVCXcjco+TkAUa/LbV6HVfWeTTXHGPNsjGsFync
jv87t9khsiaKZGGOHdJoyPpJb9xrDfr6Aeyfn2GoOReuepLNH6Ntj6I2XSh3MAMh
1ulv0nOEJAMFqLrNWsJkqta6FuPI1XRtk+48rB34qOOffcKfELopUPPSph1ch2/d
fOT3TcKVX8n1QW6/K1cgIvuT5IHOhjbAp1pNSOSPQ/hoxcjwjw+nolzVb0Xz8seU
ME5hNnspelMMfWT2o3B5yuGpjLzAFT8IPm1VJMnc+ZVnWFDpi9U6SCtWOAEpBpy9
7ugczZOuDYJ1bFszXxgEnPFPVQfheERcpcGj8/7B1PjU2NzYSEzKW4E74JzWkXlU
7niJKsrv6vpPojInZK74yLcYH3NdMCDt+LlRnMYTc1ju0VsuH5GXxXa3f6MCqJDs
PxgL3tEBAr6L5dRHE//o2a62BeLWw554wq6tSADVlMjNQz+i/Ixf+ok7wbjR0TKE
qwU+4giyLL9g38utRms0qGp80dHXbLQxBCh7Znw4/7Rvtw4jbODRLCiRTmdTvrFP
Mb5kmNqWr7WkqEOEqpaH/2Sq/3YH1+T4VQj978XyuEdiJrlmW99HCYPDxp6MIOsS
wd2IU5Q0YWsm1eTwKT8+7JGrtUA/OKNXdk9LpZG/o7O1DDJaw+Y4HjHjFN5AcY4g
UKsp6iceWfw+2tA88zWM5pbilRPSLO3E7UmFk83eV1Iq9OZbQOd6243AoXGuN7UJ
lPWOG8lLj284r4yEfbxhUiMnOAbVkF0fIvUXivD2kgxdzs/F47id8BrzPoaTjYkt
4TvWeiB5cEGbCiA4n+qpyynZBzO99IAkLW7/8R3nYzK19ZpBGSqNLkvB3PMXRO5p
iIUHQ6PvwviViiKIc2YWualXhBrSpYrrZR4+WqbV+oUfGPNeoxZsYy+Far5a1VA3
RKUEnXULe/FG2ok+mb21NFNpcCp+RUvlMMxLOVhpM9gzzvbmA9HWtLxBvWuC7KOK
DtqrjUiLB1zcPWe0p1m114K3q0pmxsDYeowOeDwtrcWAnJAQctoBMdb2lBOLyfRY
mFDJ9eXsLC6EC4XQ+U/f2FEWj3IERxLVGQe3hePe5Ak00jfMWty5T3m40tsji68z
UmhBy/PFpqFXFf0DoPTvJkELS7ATGzkk3O/LQSvDOogu3QrnOb1vbKel8sqdJ3vU
HLoAfrLoQGtylb2nuZxBivnmUxfZCvyzGOlgVYvGehjgeIh2p3Yf+n6mrgXTcjJM
+DSReazksfBl7wkWGxMForKguQwwfn17kfexPfBzaPlD0HbeQiJJPvj+7gxWhcjS
8idMjQHTycbXO7PPETNw85eWT5GaihbUcKB+DSvx8HMZf1rt+RoofFrtvfC9a0XT
xLtv5k0rkixfjxPZfmgTS2mchpaqr1av3iyKkKnh2ESdV+/j1LlJmCnE1IeAn/Aq
6UNpTqsduynffPgX064EBcMLRZ15NWQL8kslQJrbgoOac3minY2k+xcsVp6MvHSY
W0HrvQCvh9UuuCAXHd+BqSJc3dE0vNyu8BNqHaDDxqZI4ItTQX+JTnbgQFbk1Q9t
siA97UXl5jo6JBasl99MoYtThWM7oi8OS0On1HydgpKef85VQFi0+LvAJZlwlr0+
xp9BG7v5mGaan118Qf/6wtKFFFXYoXqk9zVJmme7lvkgnCNuTG4zycQ78pZ328Qe
tyGuhO4HMAjtSGfm5zf4R1jZBmcDpWYxXFDD/WlhhXzYnKcfFKufGihANe0dGnTM
TOvIQyMuw3nu+a+4+EOKbMfGhxBTiEqux/Slb4S1SFPUwygOJ+64hp3eQknfbz4k
2wL7lDKrwxf1ORhWpoHLNMWO27gBQPUbMS9hc+v8RXh1uSfMX7KTxi42KZaPW2X/
XtCkPcCaJeQ/VF3QNLK7kSBvkA2UIdirtNie86c1T338+j5PqI2ZcRWikB+8RmxF
BxARe7ThFjC3j9+8KAUjJ0Tlf7IV46hAn0o1dgSbitBhxHQyDKNP6riq1ODKTSo/
fUO1dH2SIWXlLoc8o80Ue7JBfTFcapmdE6Nk1yF57VDPS02AEk0IYMVp6Lj9Kh6D
kmpGC5GCnwYtsxC/3++myCv27UqaCRFGPrRoeyg7Y1z9JCzq6WuW6/KXs24LZ+HD
EU9gTbCXRF9v2b6d1R47lJA/u2ZJqcBugIpF8hYwwnWhkrrQAkLS7TUO18ltZSh5
LId0RnM7sx6PK4X57F53koUiKjYpqrQNEIWfUbeq3WD602qfrZgbjZgy0XZ4Trdn
MNIpo4du6TcvnFzH9MPoWvTVWLQwJdBgCBbK3G3jpBR5iB2lFWEzvGvXgdXF8pEx
1RJXPnZbicDDq+1HOAVXITifcAI5vxH5/zh97LUMmIl9W8TvlBWA2XQFPZpROtxx
hdgoKGqK6/vug+wi+5hWC25R27xXWZn1V0lt8Xwlmv0HBIFUzFzd+haz5NHWkwcE
B9pMk27YL+s+KGJ14Kt2eALx/tHQfmy6P1qXbLVBRf+KeI0DxjpCJWuDmsAoIFat
M9CRuVVdMk8wHmAwxoTS68e661hXETqCC34T+CWANDmNqkcxt8Pq8dPa/0nIuvMT
LDRuIT2LysImzH7C+fzcwdTrQ2XIjVmBuYA3RFUEgTaIK39hqIzFRUd7RQ0yCQWn
V1Ui0Ka5kZONVQuVapEWSyooSsagoaKkAtDGyIjfgse3XuukVCuiD2fyA6T1Czrl
Vn1YoRG039tYfRd9Qr+uryxM2at33p+ZY9m8lb3WzteXD4HJbyKbau3DlsNG0R9K
9DlbNfNF3TLt3JR2q6obGrDOTN9CjX5pQ14eEfFA0gq0z105AQjYVOoyCK71vM4m
tSaGeHz7OAW/tdHMWUrDRZd/H3qwnZEgLi1Dr8OTGgnVOKPtmuqxTOVdQnMKDT1I
xdqxPBNaWcPmsLd0PP7i4ZglnBhByu7pY1NBUwl+xN0KmmgaYZvBuQQ8w9t/nAl+
TGhF5So5nDhVHWkxmBiBnXKfpPZxnyKjtmAyzBQT3AJCeH8wvGYFgxkZoM2Fzmzy
IuOfpJzMfA0h44CmFbBhXBHoBm6SWlLxP74XhbjInVBYabXkDXrSmvoQu0UTWGxb
jE1kYRBc7y71rD90XSEAFiuddYcVIXg+IQmAN/yL5eNvnHJTjC3ar+Zw4Vbgaavz
Q3DkHSps0VEFx/0CAljM9/EWZTl4vd2fvcidCCwJiZ115oCqenHNb1E5tp3Zxn8F
KzgPedqHHWNYq4Jv3EfgujGtu5uxD2/yg+KN7XnPI/0A8kc3TjPYT1Y+hvov1TXW
yuwlgoSCPNAaP7BqVPG0ArOyhfhEjUsex0R5qsjk9XIKUmOkRxcl1ohFVcdsCBQs
haGktkZNzYFX7zpeGW2TnJfdMxEJy70o/QLzdM0iwIrwm9pDt/ciANBBVpq7jPOP
mkKJkM5oaULnTzmsTjn1GuFzRShNa1A1AUjkvQy4dbw7SKfMDdie96gw0oOByskF
kFl0D9z4r1AoXHeLgiUOe7J+8bhDaroJfIUZ6OH6mNLXh7TMZTXTL3YUwMs8WIKf
n8OK4dpi5x5njhj0Tcem2wLRCqk1f9r9/SJ/t4/V7iQI3c2zz0IixhD2nIBVnceP
C549UfitetBOokXjud8X22wYb261hNwJCl6DoFpjzogR4zkNzx0OeoGU1WA2ZFz7
ZQiARPhCB5klrQ/uaP8Ux78UDbjbhe49L4jQQMIdCDEOcGJ2w/LeNF0jmejZmutZ
SBAfif6bJCQGblWU1dWMuV/Q1XIBYt7qM/dI7Zh2Bx4zbVz3LgehwuXkMcWL23p/
2nwxfcoPuOLMqz+uiY0oomWWKa8gQiFKFoIrSsc708hTxdlElifp5+3kabZn1gqK
byeTDHU1Ilb6itQyCNYT/cTNigmr1GKoN8C+z7QOyOVcG7VoM0znyIJdU3pFdngL
ZavNPVxAkGuaLyZp0XzBjzK6gcVqdhyJwyMCNQIhNE/FPtFtx52G2AuFfuPEJjYb
Wkinn1JjYHetFPw2QRt9RF8tTdcI35RHWxvdlvQWWje5Z2LUJ1Se8Xie9gjsoXda
cpMbYzpygVBPvtyzAwTGASw2IIgNg766t8qaUxU8w/JxeeKiIPRIJhL+3NyRfH1f
+gFWv7pi31xh+z8YtkAM76mubX6EcBLra0dVM04vWKcTkIahwD0gHyx0GHyS06gM
5hSjCk1vqTUai1HLTXvIJTs37EqHfJemK5lX+WRDpoVyeSA6Obwrmniz0tVyApFN
n8xLUELURbXwc0aNmg1QdPZ44oFFYE4GwoGAXS4BEYRsMNxhXTq8SisfZT2bUlgG
cCe8mrbiRrNox2YcvQvhxhRMygpVrDJ9ETLa8Lve13+aiofJseKW4BJH45YVisKE
u/WY79DnNjDzdUAqcBQQcgih0aLj17eL88KiTWbh3PK26yQCKZ2NKleRVTVi/SNT
vYK9WhZqtmhlfurn6YZaThe9CRJdN/ssxEAj0+N4kXSNTCKf9jjaFik6FT2eKWWn
ZDr1nitKMDFG0aKG2XW9CF/VlM/a4NHom88/ZPSSpeAGxsSPSyXGuZfaYuDFsOE5
0wKrvrivCP2svgB8OeMO+dX5cpTuyfteQnPS3KJ6Xr4Suw8j33aF5loajEKTWtBc
K1GoiKVoHyutq+WYGxa2OLHsTF8+ZZkJRv6IWNw/0YOtzrjWP0qavvfSBcymAhva
EzYlEUqtabvCt5pKJiypApZxQBi00qpMy0Tm/il/qafrmpbiuJdzhAgYpcMZhNH8
9SylrOkFcNRoNMxrwAfey3NjsxtYmVjKAOHYCFWL+5rfrSsnJ5QqriamfPi8Cwr8
WoAGVtVrqpMwkDBNym/Dv6GE8WPcrHfRsha1OjpYQLVJmvNA75MkwNxRxjaG9ruU
MNSd8ji6wngqBYrK0GzPwnu3Yz5YDd4U7rR4xVCT0p7gHS4OrOtYUK1xoTrNWH6p
3YL8UeCEw2QcZXGgDgmhxXzp8IuZQtidloh3W8PDxL8yA++VFJc9nQWNUWmEhXlX
p8JGXtJNjnpfAUna2kmqKTlTB6HizOSSNjrELP8vYtfKOIBk3gO71VH9APWKmXMY
6xr/oQ21yBIeJ8TtFQ8J8rZ+L0GT/U5klSu5nxjqnZdwy468ERWQdsbBqCn59gZI
V9haGpC2OVXa0fIJX4hnbVdQ1q3lcHHVIVrupHvhQ2xLZXgIHVt5O1KQuiHntTa9
31N0Tuf7xBkVE1oOen3CBjIlkhkZHYQ22LoIZsUTpmptHqPJa4HGWHdPhP2fzLBX
xSZf32myB8H582s7HnLQi8LBDXV5Yp3ISNrdRJXDLR+QWuwKQzZFE+zAd34HxGjO
wTX06exL7EFRZxBk80eWmQkP6XTRY7A7wgaXVyOkgSJHyx+GqQ4X0wiWPKDG+kUx
BDE1lkWySjUdHUvZwvqj0YJpL6v6Ec7weQYUL2/k/G8GyYadxiWcTww23qqoHl1L
7ZYGBjRcH1slnEUjFGlLTiZIcKgNnDoynEleuwi+0WF9ZC/uRJdTYlJJYOjTx4/Y
WsaZaWuzAN6eWxRCYu9EwbfpeJfxyvhjX7xDFItzk/0nahIhgaQuW1LQXX8tQeoN
oyRLjfqkY9avQI5e+nUVNAGTmaVo28VIKXzxpBRBMRxMy1zhhRv6D37uyJyx5LZh
3hfleSOmoZ6LZtBY7CZc6eaW/4i/Yn2pxrnutS+3ZvBiA9rxdoI9DclpGMg2FT+T
1KW9LcWlCrd3mfeS8ZopiE1xrq2G/2lf6zRAeRiwnE0+o9eSNNxsaqaj3D3sm7t7
89DRToU2usxtVV7eUT7BazkfVnp7ssSZ0cPoR9SaTzGc3kd/80qgqhhcVnAHaJ4a
hkETSVQWX3+7H+5POe2wTUVs+hiTmolLus+tUXmLPe1bjeuW4DVe9dKlQfLCrlTi
/hV3TSaKzjuCmMmZ0isg6LFimG0JrraK2Z5ZsYFKwl833DKMaGIz65yxV0GsrpL0
yms6NWvA14qHwhlmxgyCOH7jawaF1oJKXMFQpQZNfpOdmIHvDru7IaOeXj32Pua8
YJ918NSGcitdkWfFYLI4loEOBCfCwWSdOENHelNl4kw/SJrVeuqQRNDiN+TNYT9v
CawnmnTXOByofgEM5BnhN5OasiS5iJPBt5qdkaAgcOR5XWTeVwWDYy7/Ww+zZXE0
gbjIDVh7ob8XnK6ev7FY31nqg1swpdAx/ofi5fI24H44Gz/Q+SeKe1ycvb3h+NHG
sSA/k+o4RV8BQufLhZQd2YiSeygs0bTrm1F0samSswX5aMmqNqnB49XZYSzyb3gc
S71HXzDtkrZNCxsP4Db3iRXxxk3aMd9ev7j9iNHH6u9I0wC1HoZNawwBDWUoIMHi
hYR2U/+b2L0XroxJJ6Q49FqeNMeyVSgCokneHnuw+YroUX3jEGX5aJdGyEYSnyLN
I6sVaALS2qJwFmO1uRaYMqSaNqCqLp/WBPhOBlo4f+F2Hi6hdw8SO24Yvi/Ke1iI
8Y15XcKdYNVEy5L9kgkt+vpwt92ssh5u8qC7FiqmXARQI89Kefs9/qumCGMSfFIs
/mJLYHotUW0xbjl9QIDgQZIpNntLYVaJ/67KjQnmX+t9B4asihWPsERStNhFVsAa
0+Rbtl511trZz6XvaOrAmirffGTXIdZOwb3mld4QN95A5kdzROIAG+pll3QR2uF0
ryjH2W9WB2TAKYzHJgOY4nPHZLWr3OhQzbv8HNksGZDOD+yrtNuxCTeMO1WMnYTT
Ggo68DMcb0KqIddG461x0ayFgpTXeu3TLKHoR+CPCp9MOs7O+slIf4G7W4kyXN1x
X3O0+vJM2ySn7C3RzJoFVqKgBwy00SYS1HHCL2dpAJCXgAqcyMTSNIdzElmnKBq+
JLT3LV8xDWaV8i6WbeyUReaOqfgwxy1S2psCVPU8g0uI4FS3n6bNwbxBtABUbx0K
6aR3rsQ3XlAEhF8DW65JHt2Hi0vLSqIrN3lLo0YxywxhFeS+M9U0wzQGkzmMM8NQ
2OIH/KlY5OTWFDfl4SyrhNAPeF6ZdPX1Fx8Ngrg7OnK8Um7FUygOkUgAYyy8LuST
EqNHAYC3d3dxbQgJZpGkfgjw9OECkycVEFq0qxmOyt9pbDXRUFX/Fi+Wq9MNKol5
66J70pzwV5tNFfYp7rNGzHhAnMvthSo4SpNDiJKImNL872CmkDnSs1vnh4lKmtzs
nPQkqjhJcZvVH9kFoAE5eJ4Nk5sHdnEBNT1J2EcWAsfI2aqX5t1CDqq+Egj0YUos
vAqib9wmoD+JOamw+z+GYRIbboVyLDABglTHwfYnu2qakM6unWJkbJmfCTvHI966
fDmcp1AwPyoVdz+38IyqOKq+tSgNpTwWWsGM/YXyzdv590UBNWVZeOAGnUscSZGi
LkePhz8ui+zdlPavbaxHMH1tCGdOQo+fiBltmVMExq7cjkVy+Cx9PwL9u+y7R9+4
+Rzo+3o9hN4cLTALm7Zn9AGgZWSHmwMhJmIxTiU6WeOwgA5iLy+dKkDIHaWo6LTe
sjjmz93Y7ucZSIIiK3CljYT0CuXdwI4gyeyXa2AcM8b2+wB0JbqdZV9fxVWlT0pF
Ik6dDhVusoWzERFyR0jCYMy1yEDOql2GH/quC22l3pMHwiRMk73Iv890IpEg/D78
PrnaZch89An/KcS+1CrgLyDq5JBsre5LN37UpB78+O2L/ekU1en5wACqyc/RBl9J
Soy4gJ/GWJS1uG35va+12qWC1+AoulxOL6onWPpTpss0pWpOmakrPViWw0UF+9oE
4tZee7gMF+cBaDTJXhkwbFk5+mHm5LTz+C5gByLcCEbwr9xGqn+Pm5GNz06oFExz
gmd5dpRWeK2LQnwjJ2qGR616NahzGxQ2NczICHP1jyFJp8WztGV9oPWyLoLgqqJJ
VYuz+6rGpo/OFbBmaBAt7wzruLueja1Rs/UiE6RchWCgmULXx+sPJ/Uppd/69pqa
GlL7ohDmEC9XVw4N+dLiFKJTwpuYRE9/QnQUkt64REvhz3bgJLkU0vqZIUpGf8D9
iDAlWvNq5UQpXR0/Ana9bOOi+0kV6JTVvg1cDzOSG9A5+8ucNjiYhSootYhgbyGU
x40VrKBSnSIAcSb7UzDVYS5I8BW6L/MwZAQ/0xJf00LuU20jZj//d9Ef2JZ//X6U
yuXHaBIlWfGw8SLYxvgWxgF+lW82+MeJwaO7mH6959RbZE41snf4tN5rmfw1wQ5h
4E0Mnv6ZM8JPxAByLK0DF66ayzw0KPNU3xEg4diz7oYzBYuUw3tu6Emruv58V4zc
EZIW4EGMj0pv/523iSTZlkwV4Z5QcD5PF1cSXImTq4FGkf8HS4nRvTmBYKoq4hWa
k09E8JWXmktB/X61nevfY0UWEQIlWEWkQuszT8YjIjHip2izPudVPoVw0VSD9gQd
Cz1/CB8vL5D5CkrKdM7DV7VMqqGIDHuU8z/EUjAdDp1G20IynWqb4Z5rNsVI0WHX
Qg9CLXnSs+AKLXeDNTqI6YcpGX1hrBd1ng+C8p1bVTUsWI0X7MsSGozXm8GmZONE
tDCSwslxZDcNHrS03DnG16n53ACl8/tvT15YXSTMVVaJwQMJjNSDVpcPlLBNE8gd
nqPMboKih/UkZJkHywA+ntcA5sKs22C2k7aytu2bhz4YvXQG7SM023aZndOJ74Sa
1cLeiDnHvWS293ir47msuej9rrofgODra6uWLZPfUcCk8pABzzudKfoYPClHhQWf
lMquMXf7HP3HZhdM+DpV98pewQEvFsPhqErPsPkaKTV9K1Mg0bjDPMfBPjprnVJP
AoF1+4svuLce6RnM3topqXVdgAFgkzn9nNc+EW4TPeY36TW0U1MMtetvY4AH2OKd
9KZJRBxI+rHodnKOA8pXgBIFKoONZjv3C3wejRryslhCHLrOdBQ/XZJ75zkTcRqu
FDFmNqDPF/TvqavWBY95zw/xPKJdzIU+zYK1YoP7cdsJtErjB7ajOck1MyVLiQ2G
wGQUiAilNJEkzjHHLrrJFkikb7XFMGmLRjLzTX17nSZwNQ486SP4b/FhSGpJNgSy
fwKu93cI/UcvlHR/jX4cXGB/pRMLSURjsQiAhKpC88043R8XqVnRQkOAX21gS2fQ
oX8hqKSL/ZZBcSPz9G4e3zaKz1ygovCtuVE9Avin+WmH7S0y36b/jhlnfrY23a/Z
ii5zp/4sf2k47btpVlO/I/8gRtLsnFUjplKOfCUSVTyKPKYPvJH56aVoKGzJXNBv
+Tfp7xR3KwTvUxuT4icN9iSqeiDPVa5trEUBuyQAp9sqMy54R/YSBT42NceM2rP7
mL+iac5aVKa/R4wyrKDSWiNbuboZxT+StOWIsy/HHwgxw2bP3OPm5YafAtGr02gL
wgNV7j9AH/nG05WSg9URgFkcyjBwVWtlO0nLmTlH8K9paXROhlpg0GRHxs2ej1yi
Ee4jnPQUL2cbVsE/3hp/jE6xsuy5LyNRwgpetO7W3Hlw9Tb8IW/Ixt+ECtkOO+0m
rw3m4Q68W2ttW+2iEhj+gASTdFWh82nUFj66Q2N8Ba1WuMO9X8+L9beqmsqf/1xI
1QAgwCM/zFosShRgjWpEvtePQ1xUYGNQWyKzuJa6bagzz0ecfZLEt8+TSNbh6iZs
z8aKiwaY3uwZYwUwAULLeYDrR1BoKeHRWxH8eN1x1h24dNDjctrAYO5B15RPfPHg
sD/dRWl2OKa4JhUHiKnb9DKkr3duk/hSkzgreJnUusxjyfZJLzZt6TqDWklVcfqq
CN3x+gvVv36IYjYNaV6hOPD9FjBngzfl2T8c7BrpglXs/uKWMJ+iuYFQ4rPsI0jH
qs0rDuyAZSD9+3CcYLZlOlSiAAE3AMlHgHLAVM4CIJo9X9P2dFajlGr51AzPC1jW
vxLqMZ8q805Kq6BW22UxIJ7DpyxBF6GpK/TjRrykCXDhJtXbrSMJ6jzYTmFqhZdZ
tntCbeWJ6jFtmknIhli6X8jinhXLb9GS8d35ZuBipYwhxUqTiXkEo0PJ62i8xQUK
xReTvUj3pXIvpscf0s812TlhFYiOkRAvWXffm1DPXjQKQHDJQzcsBZbvmITyhFST
bfIu652GNZlWApM+szy2OFycSrBc4b43xtF/GmXsTNUh6HfsBcjjSRjdAchd1JWn
tSeaV6ya92kS7hNWxUcia44NM8QzSQ0tJ/YSAgVzzSfZZ7xwWjashUItftrlK6dX
QIQ77qzYFjdxYFB+d0j/AVB6eRYwcl9CWfyMETGo1TSEOx1e/Vm8cBdonYhAwbEu
VbBG/4p7IRC8m7EvekSIUYAt7TkvZB+lcRK7OsygLPvp0Bymen7jrAuU1+2Ew6Ra
UwxvXk5SBB5mKUJfVrB7Qvo/Qh3H6KotO7/CIIFWJzITn9w2Goq+7/WIX0laaLGt
fEIZjpY4Fq2b6538JHCNBtN9VXM8pardPgIIbGYnbSeQbsz9b7msOCZZQwp2dPom
Jb7qdG/a7MFxtijg8Qa14TiNjRSqafpvZnJmz3U463OrwMNtvW/nZDEbwWPSjMXA
/EpRVJQEqOzS0CllkLLEQ6n4N1hQIGBYh8GgEn25RAOH434BUOr+MnSTMPZeV5E2
3qLrDwcGq/q8uLNDtBFdSpsKHIuLQxYvNRCeS422Kb/9yuWyd4J1bL6Z1qmdsTop
NAew6waGZMvbsPgSMuKcpHuFkrnrS+sQ6Lv+eYXd//+8u58U4Mp9CuQhMkT5prri
Uyqen8gIj/SQnEJKAlrXD5Pcd1/M8GVPQubmItxBTAkl/9SCoMsDvO5Q+VDoFbZO
wEKvfj5fmx0rPMzft1sLK3yHcIKkUt14qKc2o5NiAGXgUqsqDsKk9VoBOSiIL0cd
VI9hrYHJqEXyR1jb5ZJr0RIEsFRrn+iHzP+HIlxcz2ZMRixs40ylFqt8h+x3j1c/
DXr/aEzZxPsKbbqupPP5uO9XpKXCf2Qz6sSAktuo0kcxhk0bzhvNusUOwtFMmo7j
P+aWg8FTfEJRhVRc0a73czPpEdaU6Yi2dPefCf4lhSjvOV+33jmbicvJ9D1U8Cqy
TCtcGlkJLQG7+pbyrT6LXHkZj8b68J5bvyHEdxW45KPN0q/pOab7c0Yik2rXfb0t
i7uX/3HpnjF/hsSQYeM5v/r/mtFADaxOIgXRxVovDLbkRSzC/sKK7q2myqTU83lZ
y+bzCwqtuOpC2x9pdcrD+9oCLUpGs9DOEkOsI82AQtUtGVMTrmuXrF226u5HT4JQ
+Vvi72t/wvT/9cxArwsszUTBHcUhKDfXAG70ZgfoGeaBBD0/9r2le8qACaWjHD80
mx/6yk6oDkZmbgJTONP0hZmnbjp+o1k2vwGDTV/UMDopPm6uqdUhShG99nqSxrXm
Mqnr46Sc2XLZV+dzcZ4or5v6JSe4TE95SQOqEtnaWeVKq3k150LkWE9WAC+6YxHk
mUXapF2ehI2Wikl2y1wwje6A9xIEt/AMjJpT4wpYUTLQiTko4eu6x/CZdTkTzGo1
xjg53av2byTsyHqZSaHcIHKKXo0BDn0FMGDURnDzqMY+yue9f4RgvvGy6GaJvZ2X
uSfs4AJHLY9NlaGaZRlmbulXhQoT4Ot6JHbxuMZ9Fwe9QrMCl3doYjq3Eet+XCPJ
0Do86xAyoA+Sb1+xjyVWkfwQan/Is+7Ee+BtaDgdkE+Hgh0gFP0UIsKzXrWyvxQv
r7EUubnpmmwabISDGbCWXzp6j9J0gQ5UcUADQtko3CGECBqFxvYI4PKAdYl9OTav
bHFPtdvadUVx/xH/rOmWWWQ5uyeRx5tXsNUG2vcv0s9lyHsqyQFHy59dW5gVjYE4
EG/yMfmiTZymtIZBvPoV6FqC2WafcAXuspXIdBiSttaZP927heMMmPq5keOE6ASA
zDz5ECcXwegrZVzqc8kG/OjuhM3jpQvIY9L+UJylmkeXL2JxeBtPlwq7Bw9Wf7hj
eUJEr84IanpfBEw0LByyfQAMyHT77Nb2Ko0aVJqkbv9BtIM2YptksaIW9euFvgtI
zi/goqePaeftATMS0z6Ayz/NCSZsejSGvYrRrIJ/AXg/oaT0FtI/um7vrfd5xIZk
bBt5aG1uFEQZmZdfrBiLjBiHl74kGokYwWwabkreFcOeP/+WpUxE99NtXQ2rytRp
nRP6KBq7KD4cPIGA5HhxYaQozQVa0sEkb8nUHJRGdnBu3OpkboLTnaHUbLnhwJqV
4NXcZXMi+bZos266WxI+wwqh4+VPru1j+S0RQVQouw6/w8SwQu4XOQ+KQrb97ucx
EuLaaX2Rlc4sLshIMlF4lBxnJWsht7lnm+3ahpc4xsWZZZOu7ldf3x/gi+Fkvd8c
n7sTm9WWvSdhOK0ukgo3z30I/82i3innnSH3qTXuUtHWwHl+IDd3eHZZ0w4FerF/
GlnBNTUBjBkfub0hYPa1qxcQabpktcE2SvUZiKNW6LbWXKxAcNdhhzEsUm+or8Op
FOm6D/nlpqEzcPPj2KSvJK1Mg27ELV3KhQ+7fyYIwU0swdFs9egkQMq3vUOE9aaW
90Rl4rayNK9crkNKahiwzxNfHW92likmJ5D1RAAXoqmAz3mj1Veds+LynYNdLV3k
rd4wE1XkeIEKc6Pww6b+dg2f51snGolZ7syqXDBcJrnKLygPrrK1MpS3+URui7uW
1JQ00d2XssBhHR5O5Jh7kUKVomEFo8ujqNNjO8MVItR0cFR7HcV9X0q2vT/5U57W
ojot8IFVJ/+0okHJmJCHp2yARUjvcHxJCd+aJOsgPT1vp/+5x+STsdWg29lNNJpv
M19spepjo/mjml0Cqy6I+KkNnztCN0ZfIblZdu1TT01oZCETvXGe4tbE5Yxx8u9B
K4Kjp6SxgbRUOrFqj65iCgQv95feQrg8xs0omNfq7L7ZhJ2SnGI17+Ln4Cm0a7QY
+GKA0lhZDAg7Zh+LvUlBaoH1ZyrA+t6dSn/DlO+mRpRiIfGKtqQI3cAECppqQnmJ
rOC8M33rJjN8laAHIbyDuwiXue5jvEM6XjYzlsgzfPXN5AERfhuF6125kuHDiFwO
YjM3DjY6NxfseQRolTUaeb5UX2csnrOknbAE3MKRcRz6VCCrAqz+i0HjSwuGMiX4
9gEqQ0Wkda73aZHTwttaNg/PsDrPFUORt4RuTZEggxiLI29teJZQhCoQ4w09AwMP
v4jqq9QCrYQ0bEC7aB1ds4vwP0XuO9bt+PNEW2m1fInzLPtl9CB64mMVUHeUiKZ0
elqbVKcOuIfd+Q2O+n/AQgpQiRpratT2YFYxuvykJ7qDz0DyL6DEqOkvmejgQ464
LfgmACHqBREnGUv+1PxX0Ceeqgq8YCqJR8/OGahaKpOTDO+lWENTuYjoS9x6so01
4KjH24L6Dxy41Rr9d2kdTOJ+Y8x5alueeevrFeFcvl+Dmjy3TRmJQkJQT4DtA0vF
3JyvXuQXwbD9U5mlrrHSacKTWEwlYTIISMa/M/Twm2hhLM9k1+HQyqlXOXoIbKSX
IJCHRmkrppWDYcARx8KIFFM8TDlqielsR+2b6tSeoILZQnQucyRysIVmzifDSxcX
Bl4OK/SPB/O9DX9eos870iQl3Qp0l+sqN/soNuxpuQzUHtSl2Obzk4SvPCpR03Rn
RDvvV9SiW0Q5i7e28mPDs3XwJvs4pgTXMQlcWZ3mmfCZHuv/zCh7c4Y7KTKxjzuK
V3MINqrNCI4boe7GZ5M59PNrQyfy7zuFQOLRnk0OY9mRxt8dKUrTzLpVgR6V78QX
iisRkECiwovzjUmXqswAA2P8HYJJ0u0cdrQyrCyIBGA18S91iHIxz6jI51c972z3
QCwbdUqdubPW87bjbeuAA8QbKonyg4vlhIlyXmXr+cpcEwTuVBQLGuzxC8mwaPic
arMT5LxJGjGsJoRB/uXTvhZDD5Tr6Ll0qpPCNzGG7JBg8/Lfb+bagb3JR9vgukqU
+xatA/cl4ohTdg8GlxTNndr+rt3trjjLW5N4be7x7tnH62907zX1uPfcfng8mKBR
QBKksQCSlKauKWHD0/rKkOLnndyaImj5fUN3/77vvk9Q7y8V/uRiJvKzKMgDxIPw
zzPExfrhb6O/ebD3x44wCxy1IYzF0mGEh88nMPfSNpbh26mPyqMCIeY28rXgjaiP
oqaFBKpNth6soTr8r0cbALRYb7YUQyXzEKmqdV/3NFG8cv4UZ/1FlEpBMR9M6E2v
U+58LNSXcd5aRvZToe4VP87Fd+JE8AcgEXxgk8LkDC1P2qw5ML/gGsU4JE8621wa
3rC4MN7CTGj8nPjHSkTnvJXSA3oyYobYvM27NRjL3P0PMSmWyW+VUQS0W83yx9N1
jLG8H17mXrCdki6JeP5cGx1DwmyAN9OZriREecpnY4B/hHSatcMExeHvR64wPJ73
EOaqk98zSkXdDPZCAOZRbbmcYoEeujuBPMC/oAfyOIr/5xiolxUQBgQdixtnDLIi
YsUBFI+1tA0t45jPeP96lEQeFYapu08tErqKa3tNp/PH73ooRHBioQktUXVClog7
bAD2HYBraJ0HY4BbcRDavLTYrNYZ0TqX2m7RnY0Nyb3LS6LqnZn4wpHHmb/B4/tB
C1WwwVCT3TRpJBdTENGZvgQu1Kj9zDh7momPM326Cx3MNGddSdxRCMXF3Um0qRj8
MrJ5dwkwPFh2JyY60kT5vXsVMeLfTo1SOGqB8P5bzF+ZTBPS8JsOm+lmrKPUZUqj
O/fNyaMmlaVAqngraMLmQAIvrFVmWvsHgBc+LySwzkFhXberhk0kZ9K8VvnjFLWr
azPxKUBHhZ2iXk/bpUEm0HS4wTeDonwZL2bLGrrLmriuU+ZrBCqaNZ99ydf9R6cW
F2ILLt+7fZ6CpPN6jEEVum4Rc+P6U8QvoW70PXpT1XfAK3EnrblZI87rxtaDcjbZ
VzBToSudLphQr7xnOmdrkBS2gTLA+5yKxiCpj3MtSz4hEjyCP367l9tbvkXmKV5s
xyjRgIq4ZXIX9Pze+yhgcSsLRtJr29tYDxeQKtYCWgfFfauGsbXvofChyJhMWyi8
MgFDWLsGIoZY4uU3LowmPJ9fY1WngSi3Ei2zpA1t2TA4sfgoxwp1NGSmtUno3oQU
0178SrhlUNTLiUvUpkELYcgUcc8wTEEvGWPJzife9Cw4jZZeAKfnjuxI1WXijZaU
Syz1uzhCG4fiy3F4N0xTFmCEQgABVksjt1be3NrItrovZ5q12kJqfDF1H3l1AxM4
I1E5NbahhEfEZ2onaH5PUXMfVcMbaTZDzu4hjBASA7qMnMtmDJIts78xhE8iYCV3
ZbsFacZHnoeb98g0Q8MNxYqMQAEZGB62n9ymGjq9qI+hMieLNJ7YXCRnDdm0xHUw
VwG3+xfs6yeBVXEN2s+2MvfnoAdYfInUlkOG9dQ2a5jrt4KQM/KwAKF6fXi1BeVu
T4duRqpe/4iMuFQdgt8AyxHLpQe/6ruixmz+rvfhg4IBsoU3rVNw5+0ZGb+phmfQ
99XowpaRVK+Ot6ly/jZ+aWq8fIAQmoMJV6XVcJJLTyQnokiCZf+Bx9icvkGewFpj
bwILsRX3/8gywV3DfEZYTunG70KD2lnlP8FAOlfa/wYKVZr0AmP+Tpu6nwiYew+r
iYIPdC/9fIkZN2+tvH1STrg9XRPkmfRpes9Qqff924lznmOX6SYqKoGivL71BDaG
+SlEPbwtBydKwXHjHjRpL1ZFQZrl3VMu+qYD2RcxeOT4tjXptIzAQXijJ+Ltn0zd
dBeFk+zyP6f6Fd3oLNhqR8wXj+Vnrj0xQtw7wXTV0D2N5Yj2RGYHVP+PqzKUhCg0
jVkXUh/zD0lubwAnAvc0VtM6az+UJaaRR6tmGo7dFKFH/5VGv5VEjvWR1tjrQcbG
/nGuNMbCF/XW+F2gpKyMHRehZoXmcHykVKTRN6AzbYuTFPORzUqArTRvVcwUGB4t
D1kFKEiZsGWJwhIUXQc7Hi4uPcPaYaJ0BFynBiK+1LIOrBC89cO48rei8f6OcIpb
5ZNlAQJ+t2s8gPnmkmudix2g/TdJyWaXYYpNAMzPoRlDHw4LUgT1znn4f9LEHyft
dNTK++UIz3YH+qDPs8iRx1wc4pLww/j6fP7DARxyXJFZ7fZHIlr37R6fM1ofylNd
mBz/zp0nvT99Y27ENo22jZicoJO8D1v/Fzfa8zm9piTJkGKKBhAYRa/cGrLVdSkE
QPcd8cyKwP12OuC0L6vc2DOMdxElzNSr7bv9wXhpCnz2QOUTfYCD234BdfxS+sl4
2gKnsEGP+IFdHkTfZi15kV0d3MUpRxWyJ2Y2NNTr9kBq1vdNFA4TuBBouCLSdPq+
CM14hTFyPQTOBp1VUT1M5yzk7cAaaj475w/DPrzSyF2d5KRqaI+tigU8bc4UkbVb
DJwYK6jLjW2fNvq5rhyH6uwXD8PojX1FV4fUz91ofY+IHuO41DfyM5XCAWM9N1cp
NbcPl7HM1BHd84UnLQEx76erAJBvR+gV/2ML0hU77Tc89PO6HbIPs6JQdcc3UGq4
rFouX7WfzwTMIpOf8oH/Kk3aYXfiCzHha6t/jR9T2pP5r7YkrNO4LsLwDVQJ+lRL
KM0TVTuLasimiqDEB4+0+OXsrMujwV4i1ujmAp3hmjgAgWDgcgwQI3/cuzw3LN0l
xmBSW3kTfUN6QOSW86Bh4pdDKi+3abT7HCUE8Ce9IndSfZNdjDwHMkbpQNy4ZIoM
FduIQDA1bJKBmDEj6C/gwExKSxGbnZKXnVbACyV2/chRpfaAoxz+qMXuk53Nk7IE
qEMNlydpiPTonaf7yTfSFgo9NataBIay6CbJ/zAPVh4vXtnnlhCcig/fGI9syIJE
deUUc7G7vbQBEo4x10ZuIvN+4Ix8iYA39r2IfLZFYoJUkTF5R5oBZqwGKXMQIEei
E+3JCvLFLlu732Y7LHsc5LINzaZgUq+oSdg+5h3zXsQ60rJ/pHDaOIrbem1Ib2IZ
t8G5W3bNytXPb3JrZqMWfXEYPzrD5m9e4wHSvOQWwAda075cEkEyEiWFxFvBC0Bt
4+MNBpe+o4EJH22AEZeU3q12OCihbzYUENDKN3QLWJZLJ0LsJpC/BI5auX/RhBMW
5Yv299YQs62svA9FnpQSIoPuMLF/V2uAj0O7Z1ZoUKW/zlGbAQo6Df1wpgd0YXtP
ajQDUE4qPxRo6x9BCkXV8XfbpW4hmRfIRQ9VLic1ObxL2TaAnWACz2SVLGMPbEc2
JK4H1zcBeTkeNS3RPViz0K3h+zuaLeGdWFcPnHzErOmEuG8BzTFPfmAfFx9vO9il
4RmqQxo8U3Xwhk0ysgsQ4M3JynGI0yY2Y2ZIv+RnnDKzad0rFGLVp76oxR7kTXF4
H4t8HEsSLv/9mXxZKTZnRwNeaPycTbnING7UcStiuuwlZg1w1ojuTLzVL17TtSWw
gq0VxWQjPsZzdj+0qmvK/oKE/aK8CLfXZN3xRNZq8sXlJHD5hLd6IN2oAn7xvihs
QlscqoNbfkdBOUNBK64sjzIsKqWUlxI9iC+jQTITfd8xOnrPo4AHHpnHEVOlXrau
B6lxPuyJ9T0Ph/UFnDMjtotikfb84ds1hxt0/Un7wUFCgJCXhv7m+bnxSJuDwSEf
M01aXOlHn92yK8hOSd4lzO979L6Eq0EE955cCw7i2cAr9vryJ8W4o8D4oXiKcOdq
pdPMVKnrgpqbEMUKpwPBp4S+EAWYPfTeWdYstVJK9JQiocfdOQJUuIZ9DxxSaqTR
tXxQ7TfOGX6x4HdP2EYjUgZfzGATigjkKSA44RJGIRHnOSACo4W4+q+hkjg+W0pg
QFRZ4/7h6J0yi4Pue82FJdpla8Im9FwH4nyD3UhTorZMiw7dt2Egl3YSJDMXQ5UH
OS7ABqaFErBfLvWO/DyTQJblUdGmdBi1HgcI9tCvGhFvOGKcp0+1HprGUDCCLCkz
9jZwaulm8fgvSfhOw4QY2MZJcYowZXro+cC9/qv5HjzPJqLX12H4LAbDQTul8Fgg
9X983eUbd75429qqHwg1IR5vMb92Tm77VOW2ITQ53GLqboYy2gM0uoz2BlaFPZo8
XWFlDb4CfKWjAasWQjk7rDEKWqjAzt0ieq6f9jaTLXdlkvxw6r9Y7YiMvM0zwbds
Ai9U//zumsy6SxsS1VmXNEdb116D+iUiqvX/jY6q5V0vlizZl2WQ7msc9pkHFRml
aZFbTDZoTI2mJWKvznZp2GFuRNEy0x1x+97E9/mmcb1VzvFpsDTILERaT6+LDxEY
jp4hc4ua7hSZ1VWeRB65VV5KdDPEE1t5/Xv5Nqw5w2fleWUrhKFzPG6HTsekRfmv
UzcIHx3z47GF+WCgWOW98sSZsIp6GoKfXXjYG9mlcEb4QQGz9+xowU23QILrplNm
E6xfxhGoYgeRhWDyqFiboA+M1Ck9ngdCsSz01mgKzg9Yky/n2YntJDzgBRSo0BRE
WhXue0c+V1c/mXu+R865ElZ0jdVUqU41o+qoLCwgucK+2mRHkwQeMfiYj6gzEzHd
XhtT0/O0ro35bV45UNfbeufV2prnADDIBCAPWaB5dUC/WqxTTmg8xqHVK2+TBsF2
2YnJ5OKPfFnmqjXpCFJKVUWR5/cFbYJuMyUG59GoG5Ba2mi8fNfvCf/Emg/gt7bp
zi4GihZf3qf/QRfPOm+UuHfoixT4PDEpjj0Fn/1FE5it9oB2daCiuWVisVxkhECP
JSvR1FysEQhpro+F+Ktclu4upfIxEJLtXa/8rfeZAHdYN3e6gWp2PkWXkwSAMJf8
PEUaOkK+BIKHzLRvx8cdQmdtWVmg5ZS3VdiSwJ+SVPvqG3w8yawxROVMndyoLmNS
vsWB4NbARva3/XFsXw17P1G6qrWzyMn0XK2vh74EVhGYaM/AyUNgTvbywwKhoauG
Jj2A6yQHHbJHqDUBkps4fs3NFYFxaGY3QiDT4L1hnJA46hT/X2M3Am/c8bG15RjZ
0zpFEb6Pno2vRHYR+h8J3cZSr53umD2FkFrRK6Wk7hsgnPTnwO6P/EHcflE0/ZrM
Ciktx4ccFD9l2r1SWhgyCIVUC8/tw6U4RVeHU2EFjrCCDd8AnfPdQESANUOvpuE4
wNokWbs+e25o6lg8i0IDmYWJysKbzPEQ3y016sQcBNBhyZGiz3zWq1Wjx3Nycepr
m+iEZxH0gBhzvMsCI3BnS+Sh2NHJ6ndVxWQKwJB0wJsVStGYK+KHZfBWHFsSjqPK
zxob/87bAXDnXloJ+Ji/SgmBugYsW8/rt5dCdZm9rQbYViDUD7JUsN/U4+0ANEev
hEG+91fB6RngoMXHQbRFCrFd2zFdNU4YzxXPsIJyQg7cT7xMjqB8onMKPhSBBGFJ
u4ix5QLZQIOp4C8GkQ++Z1YvH6dYqFpOXIOrNHCJ/uN33n7nU9C0+4RTIDG55M2s
+sepw1zIjIusg1PEoVv8/GiFUFo6BGrBJUbe02gAuthynJ/b00nJccNHSPo1TYYI
SIfvVPe0R9WrqFEvulANRZBX83jkBbn7+1hGzvZlxY46PuoJc0HdsL1OeLU/7BGe
GBeXWGIJEcE/l3sNeEeoF4l/xbCSdTg+ITs426TcbvvAeeb3GPyDx+N3XrHV2DZW
9e93/hU845QQR6FZub71nFOxiczhyZQ0k1L0un9F2vr7nU8NqqbzQ5jzfW8mNpRM
txUE3WnavRxKG+6hbyx92JiQfiFfK5bIKz6wBBBdltBGnDAM2P+RAc1XTCJMQwUw
Twexz7CdfrB60f+pHhjtL46NIfR2sx3n42YqFkhMa/65/K//otq3iQYK1YmU7R5J
StUJ62EAa3MtO9MxH/EguyeRAN6iiPuPdYmdVOmbRGyS455QVOdWjDsILl1kAZNb
p9xztit7crZedfZNnTfQX2/NxIayFBpcPeCE+pXIWe6lcrKPuRJhTrQo0FqWtij7
rftc3WHg5g5r+yD6F7fah6Cvvbq6JdTLLKOglbbfXEnmg2Qp3cOgFEH1Fmk3gYOA
vFNbIWixoSo1M2cGXefEJfnYets/wzolgiOoYxRkLbH44EMh2RhidSb/85X/G9IA
o2xB2dRDgfaB22VaZ8PnjLO4kdk7nnTeoh+hTBkCF1IW5upScYhK1mtp4MdIgilZ
KkvgCjmS50otK+Aw9Xys17EYDX3QCJ0bBZt+3dBmWyIM57Ro5cRosSKvlEErO0kw
waxr5f2i73z2QTZYNHcA1jpd1JId+nZ1j5IF7TFXWxzU8f/oX24E+XgqBO2OcJmK
V54uHeK+CMi3dW2BPIa0qResamdTLBkLZJYzv8Ke9u0hQtxmmsCnNj8i9w/qAphC
5Mt0Uu4yYHXBn7x4EB0H2JMO/eD8roZG8o6GiATcY1ZYlf0+cFPDNybLSDLEIL3R
QnF68vBlCznJPqFoixtEfDzEt5Z+iV5dXtu1Y0NFUxfaLE25BKRzX3yyRNS3NSK9
MTSO1GhAarPQSG37s9Unu5kHMG7I2l/h81mqBr9hdO1LJjmqtjts0CAm84nZ4oRN
RBaJge+EHblmMtn6C+jt3QGuIgdJoXTPLd0X4nleR7+85leG/8P/lP7RmjOi4mjS
ptUlLi1y90tfdgoECoO1uYCO7cGThRTkpRn9R7UB6Dn9OVDN2ngy7ZhtLCWq/7YO
K6Gjjiq/T88Ni6NKEorq4Fp5vvmtJ09e7NmkTlIHYuhXqSEaatPFBWj3WfClL9NG
XwLpH8OB+qMpO4VjV7mTRJ2nLqUSCerqCfNKmIzpXqqz9Djrcu+oqxBGu6sStEg+
b5IAVpDSWI4SJ80mawRZkDanXcWNG/bpsKTH7C4+wEUn0hGyDTTM0VPqbEd9FIdU
jWnqnNEmIObHSwjXEj7jRFiB8zmGaUwLaudwUYWp6vdIrChkXOjOGHc8na/7pXyf
KBENQFb52XO7OYFD/l8UFxPEebb72gzrMOUPTGq4YnlJ5VP6DDZM8FzkPdGCOuf0
8ePpinzVB3JSlwGrdfHx6N/xY8cpBuPqOz43rwuYC61WJDuyPvKVNzMNt/nwor8f
pFMaFToIyLuXaXdYDoqEDjVTAmFamP+pArzpJgT2NhyT79avEU4dnzoULYWZZCaS
+uE6vkjHwHmDM0unUy+LfVFJUM67Qvj1U4W8JS7UeuZIapHBW1J2AkGZ0R+GtaP2
6pIGrF5Jks0+EPN0h9bfuXF3qQxaSKtYRKl104xB/jPcE1ZYumcRvL2QkRt9zcIE
mF9IjKhvR2SIewD0bsahKYUO3e420M35hPxtMoVzHKtl8d5rATUrgorl/k1/CAFY
IZacY7QSIHhNNXFPBKF0krNn8haz7R/nYCLzfET5C4mUdhHEFvkkvxP+hZHpvm1M
oLafuJWISDGE6DKvsZXHSRhnXxQW80CJf2bSwW8xWCN7xrMzgvTgg+CrUJ3/+o/c
G1FZPz0M2YoOeTNI9Y/TO2T6MV88z0/9gm8gVtRpaHhgASE4UbQSerW0Yj8nVJXp
YliwnZN5Mm/2elvT5R8BDzdoNx4KQuzUPSYaMtdtvD76SKCq1hTNLmiiOt1qL9od
8Q/Uz2JSiAZ7e4AeU5xVowaKf1hAICYsImivEx4jeLy1GzmRdi5wfa2a5FRPQRWi
2oyvYucbMF3CHX4G5ktXwJldAYh42THY+MqssWZKe2/2oHKwADyhJmqbQejvPWWO
TM1sPDXYM4PGrp2YTqyvQF9xADBgizaUxlJK0vu0h7iKEbROz/0QLWRjlmRsb2HC
x9UkaRaWoFcvXPTa4+ioBOTzYarhzfATgNGbW6TuaOiZ1qpH8T7zbijzNBD9q5ON
awpmS7iF0C+nuc3Y/BdE5MlodYHdHkMrfZa/Mb0Phb7GyZDhJlO4MlbRrcQy0ZUS
dt3TpPabUUEGiTyy339E3wWjESzK1HwFeTEYMih2p7fzJkn129GMM1/kB2Q12kQ7
SYQLT6U/7VcByXMxmShj6560quFSdgCKWG1jdktN/7Kc6hOGrHWqxxtFnKEtwMkH
HelEJ43cY8KcpHtxczaXX8Nup+lwBcORZb9/BrWtU0GnImI/WMwWw+VXwBDmK3yP
+NHLtKaaMoq5QjOly7jkle/L7EtgwPB+xK/7tPyadupu60JpomNfvlaAsUl1nlm9
oRRmPvxLqOZhIabU+HlWQ8R6WgnuzjBF7Pyw8PicAag5T6iWRFRppLv53zyX5WHP
ha8gpQj8ux1mh0Ig5ecvHXW3tS2JFbuywIfls8JBo0FL/wZODgClNgECsycadkCO
0VwIlPula8vih0+uTdG4cBzsBiF0O8h74bquFmct578hLarBDB9z13usy+qpYqnJ
kETZX+C04yRKdlDgY7Fmfu8N7u7bu7dMCfew7bf1Pu0LOhddFx1WEQNrnfajEu+/
BEV1JqywZUbtfXchsBQmOm15k5TxlQIX38EMSmndpZbR/+gMEZR0/aP0codERdKq
I//O9hRlnTfCkPAaVI7JkKaDKvqoNpMeMEYDxWCkfZPOvj63Wm5CQcGg3/E53Gkn
3y/odH8WsqQQKYEwYDbBP+5nYtpjp+JbXzkmDCpfv6CuR4BB1Nufdg8NlpleAljn
v87J460dbV36DrxZagYUzdzT8rRV5zH2fPGziiRodVZrRiwvLz3eRjW855OAaUoh
BAXndivQxu1JojlZ8xBL+UBBoGyId1XfBcmBxg+o0zmu1ZP0bT2iGV65zZNzTF0q
UoiOqL4Y90Wm2CcWJBfsmoxNpMbXHc3i9Om+l3ZIyw0YEPy7hJFrQ5nEqhti3dfw
nCqv2k+UutCjdpfdGnp2VlYEGE1pEUaLA2JomkYH/beAT9gBHYxwJDz5oxCvvbSw
5+rJ8V/I14D6mqxjbYgUJN3duRlquvHXSgFOaxWNOD0=
//pragma protect end_data_block
//pragma protect digest_block
KEx4TdYP1ZGE3W664AmRk1hOPSA=
//pragma protect end_digest_block
//pragma protect end_protected
