//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6qrQ706F9xUzcym1wTo/ch81VQpHwWwa051LOh8mSgmR+LmiDu9MEF31gIJpviAv
WJVdhldR2BqRvjHLZwXokNREeNpMxhrsgJJ+NXSmS9LAZvuQ8PN036ErW2afAQ5T
VAu0sbjXWcnbeD+OoQereubnqF38hQDyYLIMtQKe9MR1EAPH0rKBFw==
//pragma protect end_key_block
//pragma protect digest_block
wnKPGCU7sE/Sx3h4E4k36UB/iOQ=
//pragma protect end_digest_block
//pragma protect data_block
JsJbmExsqnal6E443WeQiPuV/tuGyEkTzoFYIUBTiIWKPXEElH4jCvS3dEVt/zrJ
TBS5VYVpFfWNvtBkgerqxi1mmcUNKudmSQ0GwlAYXpBKhB/xjefQo1TT7xhCuQ9E
jgmuJ2T7SXRY0vGTENaHwX7rqEj2GSV14jZ9wNFhQ7wq7kQjoifZhL6cp0vG8uh/
/2k+OuM9HG6zGxSwU4Ss7E0Oxi6TgoDI4Ywpx5j8fdCQOkYm2QD7D9Y2u3v8s+qm
T7sabFzsnhkrFRysMN7H7A6wC8kom15zIHWJtLlB3YbzJ50XC4/jvDPmbg6nS8Zq
WWZlUwdFjozoeOA4/MIvAiE3cK3LV7v2MkCcApcsAvbLfxj7zI9QMNDI/0bhyQAu
6vC6QSr4h+IQsjBx4pdlOdUQnpKdAeGIJXausdDoaiw0AeGGJCwqgs/Hb/PtvqgP
Z0cFLMf6w+aUXFOxY7k4yNg9Uzke5f01fCqNgcRR8slmcC16DI1RziiFvP7ZsW3I
mK3uP2E139BH6FnUIjFXklY9BVxojS6vTpMLcprpDH8ph6BE+VINmbCEQ2LMqMch
FG5IZwGajWsymCCCuHz9+pVPFUZkvycqK2I604bql0tzqFWj7dHmXC7SrlzpQtPm
oookrmdLOJUBWmFRZLBHQvEplZYkX5Goz5AcHpe9w40hhwBAhwNIi8TeDyoBnWPJ
tVvq1z7iRbZ6ckGwaI4GfCkF1hRHAisBB3z9UruGBTOM5nK25X0lin3UAUoXx4d0
pPwb946/YD5GTQHkSM0+a7+ZjWSwCbp2yRyJKHZOViWWjhIf5L+tYYy+anNOa2gV
epNw5zJNC2CRIhSaEp7DlOFb6pP0CDzxoENmaHaO1xLRk8AsQWGyik7LK+Owoi0J
m1M4RmMwkR0p+0T6lEgl5v6/FpU7bIze6TCDsURmfzEGCgRBlgJqq5X97ZmuceoF
m/leYp4NKOeEDAG2zCxoCY3PaF7JebU0xkviTDms1RcFxpeYJL/zZhHYXNes1uWt
xT4OSmpmwIoCsfeooSxOkHnMok3mVQrWi78ir/M7If76K608XUBJqeApIzOedTHJ
zdeBAd3YfhgNfaR5iaxmzOUzYhYz6XRnn7kEHaW3Y8bR2goeNDMBXN5jvK1GzcSe
pniFiNhiW+w+LL8cyViw+MtgwQw+sMvaPggpfAj7oQtnn3fGKOOSP4E872ndBTcc
BmGlzLcNnAzMLm4vHjkEZ0g5p6r3i3C2X8Ts1XwQePGMc3xwgni0RT5GhVnnhCRW
u/z6OPC/v3V4nJD6+MZCmvAzwLjBA2I8DN7E+2xE6zSKvfD7qfp83GNXmzf0KAv9
FXRRXxQ1eCOsMfZ4pBWv/DUAb35JUFjKf94SNLzaAxYes8TFjAMIscpjkOR0DAjJ
YWDVUe5+ntTKs/CRMzymhkjEofwev4vlOo/yzt03fplGyz7XYMgVWRMsVREW/VVV
d3DQGBc2p0UxHSUi6CJOh9qq/hk56ZV9K1oVY/th4a63k9M2MlqLaJ9hcgr/eCh7
A1Vuiwgrl4VOwHLk/OM3eOSBnQFTV31HBbB2azfnEWhH7LMnR39um7yfwqjeZEOx
aBcbNNIH+dFbDljBMGCXPRc2BcPwW5WBTQK0jYtrnATpfD0mEux1M6MYBGyIerhd
PeHgXvK1xw047jnJpVrbbyRwV1o8UclzijFw8OdlSNurGOwAFrKI5yUcFjQeEE2C
p0u1Oj4mPvF61eH+OJC5WmlhDaQ7HySnWj41FDWF0tlzv6xbCWe/zpPyNWLEVOgm
FaUSbioP/ZK0lN2qs+/ntP7Ck2GYVcUvzUQfyyt0APT+gWGlltbHS+iQ+iy3eLak
fu2Bs4F2HAz1Sv6I1tKzedTspY8Nu+Z9d5W8JuzCIvDcAHBAb6hsnY7+bSUdOxKR
ET7LBSRKaFzCrdmZsdonKS2/oTijpQTtwhuB2N9SB+H3GsMJY6lWo4W0DKooUcCg
yMQCA4bNWdU874O0PTvpyl8/TpW6xpZ+b7Kb8TYPc7pLkj4fqffWqsm0gRNstMw6
Z43BKZqQYG9219A1q7UZ5FJOIXDl6KY5rUEUyq7tsrRQHs+9uLXLF8bkYXvMHDz3
rdtirMmFqA3hCreQ2ivBvogtKBbm9mYZMbwydzDqF41Y6LgNnenWSnckF0wiTf1o
xvggooWc2a0PrrmP+R0MIrxvpji/8mUVj+or1L9/4Ykoj2VEuis6ApTeE8GmXzPe
v2oM3dkP1r7vpQ5Be06s7W6jsJlhKgwsZ5vtkpcx807iQWd3SxAYpFWAkALB6AVC
bJFV99/Fruho+x2cK8gVnuYCwCFPRqd2HdZpJ8UGX80sOV+EGtu1Mc8AehJjlVGP
Cqb20o+czoNTu6yPOt/Ae+0F3iStIsV+wR8sskDvbWQg+Z+X/35uSKZoHLTFdMfA
eGtvktofhN1fDfITnKS3eoWQfRSHvHYp/s9BZkKjXxjYiicw/HdQVsNM5TIAiwbS
1tgD/aAdjf4Wnqod9BGQWdyT8tMsYokW5b+UapxzV66ldAEyIRhvbaNZP42mo1ny
2X8JIV2Y6FA0XulkkoYbOsLI74jOk8m6RIgqejcaUUjNgpPUE5nFvLJv3zrOeFBv
dZJ6fBAP1VYRoZ63U5y6lodIjv3mTN+IrqDvInQLFZiYHGZ1cgah5Hb1zArMRgjZ
G+EKAq0b8Xa3OFOzDJgX5PFCDq0cUUEAV/WnUFklNY6Ym0EBIVjte39S38QTnsPN
Olv4dEY0ou62A0n0pV2L49tCRd9/5nPlUBxK/jxGUCCqmIpRt7nmxxReygsgQA8Q
CD7ItJ1prAW0IvOHLRtH25u087M2EAqX6aUk+kJNy19OEkAEUQxHE0d8Hf19bpwF
Vyj/gxGrxRDXTnN32h3qFENl2H2LRSDlTN/ZrsjKyt5l38eCTu6fM2q9hzEa5e34
9xGe3ZZIzMLFJ5IioIjrq9FSCtp92+XZBvs67JP/4m7KzNgs4U4T+0OPiE/uZ3QL
cNsnaKFofLT9KiwQwP13OFwoJN6AcYcgl7vXDva/FnaWaGwv6c2cAMLhRQE+03Yn
OjqAnGI42f8EFl+W0DWV+rsuu9RP/vmowrY+Folef68sXn4EqyRmA+IEZ0UMeln4
P0267G1jA60VJNLXkIlmASptUyaPzM+H0rBcNvAIc7Nwh1VRgSUFrroPKT4GBDc2
pp9JQwAQFS+DRnDHedsNrKPLjHHQRSDRAlsDNM7llKwWWDGasCniLelRdgMPgN1R
oa8JoWcBnRSmY55HLxMfmqs593zjkjH2zQlCgxpWb0dlj0r+FnySxlwmzLQfyZeA
3rIvKy5me+jzN8vfdfK8gtwHln5YMvlC3kkVRD7zSsiyApOgu1RuLbDRdKU1XIrf
RvB/juo1/aOA+0xbR13YNJ2ld68Lu+JrDjfAAgj3JPyTxTlyISQw6cj4sCwyilZi
bHlsKUhvtlSdhHYDu+YIN8u0O69pj7Lmwe9/AvBcBOQ17b2pKgyjRwlWIYLNb58V
hoIjg4Vpb2EG2SJeTNQZxpkBgz8npHplt0lZAlT+mO9gP6wQP0G+IAeBP0O1/KIY
rm32lHMbI/9xuS548MMwoL6ndneBXdqSlu1u36xatrUwZE9fW799jbO/YF6R3z2k
S4IBLz0jfv83/FWGkl+V7Uyu8JrxpkrcqQJC/HaQklzflljHZfQOgf71H4n5ANVR
GJwoKK2ZxffITTlxuHKJUn3GsdFSY9mXXbGKuL2Fqsu9ZCIDpFTL4Gr6DivUbtUc
Pj8OuCAynJvu40QrYFG8AggEk81oMSNjMduIjIzbH/LrZqDTT1rkWE+TzvjVG3BS
ODQT0TZ9PeV3Vk7B8lzkKzXuoBGm5oOoDG7FBAUeT1g0wYg0PBS0U30BgmxhaZRM
ox4CtoDHtA46EAFp2JL9+jpwB3u9RksPDzDxkowWyQbtu9Lfn3jfmghUBj0pXuBG
+bkL97PERi3jdOdJ2QpCyH1yrPhx4EptMhCntB9WqHuEwA/K1bhXA1tpfXtzpVfg
BKNO+nnHvuvD2JS4lG/HKE6rQbov+Bu9JxxNJiRP6nJEJ4jkzcygTSBuEirwWybG
ocUj6RFHalZDH0h5nS6AXwll4//dXoHAKtdgCJN/IercQy683a5ROiiIqVP5o29E
dmUkquilgy0j6PjsVb4ycOvpKkzavIIePlnh4em6kwzHYGjRGonQFS4hNjD1F5Ip
8Mnwj8pMlmqYBvLn+IN18YqXmjND5iO44o5JD2TLG/hF5EMvnT37W0cONSkXoU4D
jM4EhPLon6xGe/fkBpGVRscNPcjA6kGpjyXP78Z0x2UyB7fZWPOXmbeH3k/1F+pn
BZ2H3qHVYamryMS/8tciVPdzrYQX7+OZyPKIljA07Nzt0aTxi7eMRTYTCsclcB99
n8eoYT65cI7gw5A8g+nfLC46iXd63+PhT2SVSIBgyAK1f+5xezeTtJ6tsNdmlMHg
xTsbwtjh04/HR5bRDMTO4+s98U8PstF1qTf/NtmYqGAgh6n5bpE7VHFjEWJmmpZc
zj+C5tHOqvtfTjHLRDkSwuY9zTi55coDGvPtAmAYiJmRaNqJxTHULv9/EGW7Z+TP
67zdF+od4Ci2yeFfB4UVu99pRXUTacOu7LaSNvm9McXPjexAH7gf8m/wL+xie+vG
ydoyf2lIjc3Z8owissPS6uJT2+20xXPGRPRNdbtUG0A/AFMByJ6WTNk7L2z95JAM
iNCPtmVtYOp+pywea0OwSp/tdhALK9LDspvMnckxsqt4FNlTP8GrpQx5DQ6wzT/K
dYlxJvgWmiKbjx6L/FottIZVT7W/xK3OG0+5LmPdPPm+UMA6DXZDs64ukVHsiwac
4EAKKuQVRTI69Ivk2T3wYvwaFF7OjVNelm17GIC2Ab5eOBYeJE/++oXQkWc82pxa
tYcgB/hYlWrTcvAGI55sxBPgaEbW6LmifAOB17a6QyeJt1E0eGL1rq5yVwEZFQG1
uBB7UILxQWPANGt+kqffHO4MNNRiom8Do25nAEgCG6kwJjVk1e2C1eFT9A3ob0f/
dTYgcPjoFp46Ksc7/H7LhDyO69vz5UCmYi4JbjpynmxBJqSkymHmWL0nZAk0eA5g
i1Is2Fje9CLyOP8CUPZEZSfSEvT6D6PAXMDLKFbWfh0zalWBGR7XBsjCtiFNp8mQ
VWP+4S+QxzZSDsfBUyiUDMvEwxYP+Y7N4QODekG9qfr4XednOFCwNadpNj0Fl5pX
DfAJaxy0c6E33ta7kFcuoyGhVuYI4CqivKDuwcL2cwBZt6of9jSlZm2uF1YT+/08
whMS6w3P6IcqCKUbJGHezvUk/jI3Hs4kq83lxYr1+z4jWfcshHwMNbn4gvYO/fqX
O3eftXlUPtzIZSeviVCUYH/h+5xNByrjG4wc21zry8dg1SOiOWFpzpct2kwAdLAf
rxgHMw0uZ2vLnOfDQugROJhCwi4Hv8JoRS2lkY8Ahuy8JJJhH2PuUyGi9V5A4Xdb
lTkUcyL9gskZ/Hk0DdvSvZUFJ4MR9r0gQTcjJTs6xWxlCOl04wVNRvttkf3vnNc1
c1CVwVTKYrPdNZB0Ji+QFpA0CYV+wnXoFNm1ZboQZT2pCiG2YHKuE0oKNK1OsTX8
oaK1RGaChx4N6czt3MfziIveFnD8ctM0CI3a4wL3WFIC5ZWixGPZ6Td188ME5815
6wznfSj6GcT6RenaUbcr7LzW/aLoud3IU8u/QdjtlRUDjLKX+FttIRGMbLFyVy7Q
YhD0Jatm/TOjNaMyHFvW5R0/Ug3V3K0iSt65aL60oSDY64U/uVs5vREz/rFXMz9Y
UZKGsu7Vx0RLcEDmeCUL3aRskTwMBstdVRejDWfDSj6JQk15dAco/Km3eKarxEyh
hdKEwdsaVVlUiX5FcQBbnLBAWtMLE8iuXKzET+bRhhdqX2KtrfPlZ4TNf4qQ4R2w
VuR/Hrng1+2pQBl3Fd9BQz198NfSyIofbSNhAPit1uIwCGzrvH6w9m9QxUdErJ8b
9kdRiH6oIBrhknahgNU01IsmGGt/0iKbtbxr5tUzvgz89bD4TlQWpJc9maUY3qDk
Eii53vRw1I/hbPACEqfwJClLtAs7dwXGXX2iYwwA0NLwK1TXUMkd8fCggaFLa+vO
x/9bF6WMlZmg8ZQipLj0Z7FJS6tglI4B6gix/FmOfFjZSeGvFSv2YpSagcUfpNm+
MqrI1/7SE+k9xPLNYHkNWTPfIsr62Fw1fUiREGtAWVS2clP5FDDOF3ah6OEozuhw
yH2LZ01iZAUWsNk9rf4dmAY0lqIKR4JDUDTQ2KuCdXQ5O0+sPnBdNXnKCEDa4cl1
y8YKz+t8O1omYsIGk18cjUxfch4YknLX0wdrXIfp4Mp+mmSq/jxEsGb5X+7sjA9e
zDj1jNrHDnKIhRslLblzWRVZcLdvpygENrsN/H7coPXY0YWdU1UmiESUCBn2TtV3
fLGGaNndFBknFoVBQnERZ/ad/i9GVn/BMcHLVUW7L2dCQoPbgeusrVj6m9XAKsZc
FMG9oABhCMdxvWmCdRTAnXtN37Qpn5kWKEEqMMifK7XGzZWD7C8kSIAXhbxHAn06
Xnzy1reUQb35LgjphMU0Qmrs9ZgpVDrv8c6UXlDuN+xUJ2zszQ9XlSebF5A5/g0n
AFNtIMyFr5XZlwofmna4Ezq8pWTmsoP9FNDd6PqxUfrwP9/IItoqcNkAUSkFQqAj
MfV0QC+zP8K71gJfbd1nWY53PGqR+h0Z7vTNuNx4hh3j9JsKHUFwySYNl10YQC/n
Qdxpbejmuvx8EweR5jSHlcar1fH7fQ5kvnrCjXDGO8BE9Hc2KmsAtDIcoTFoQEeD
18/QLicBUiWi3gJXolU2hOnPkW6rH+S+vAHF4qIS9QjPUJqDwU8oEcC3tRUC27Sp
vd63hMr2qyiJMTH6Zfr7u3JI4utCVBAQy+tIHyR3nqxXb5JvJPiXgzI8GUqX3uZL
Q+qDVAFp2gymEXptiqPLxrqVLNIbseV+sZ1gQSWzT85IK56dIKwApGRSNYtpCOQY
oYq509LdjXcsjStVD4uLKK3rorLXc7JIuWFZP9kPZCbr2oUh+8AkUYkZZc7GK4PF
C9fh0pZ2p1gj05EzLnQtKGb2ZOvntg0f2CZgM8j1SD1j915Tb53y4WxtU1lWXXO6
26FD9y2EHDCFhRWOdEkI2aycXAQqE5d/LgTI9gd9xxxi62yxN6Mvadcyg7duTeLi
IC0+5OYRrEjHPvOqi/XHUfgYVzu3O0Ay+kSxfa16//f5itpt9s4m18J6JuxaRk0f
8FrimmUppw0XRdyZ+3B2FhcolhaCAoNxoe0mqOksu9oGchWuvBiY2608ge3O1P/p
1lC4tIblaNkpsPrFWrdEdgIl0msMzZXyPMuoo6l6Up+o3BlJWeme7JBWXgcLw6Uj
Ua5WKswSBfAA2EcP8t8mQO8dpyO97JGExcrPqa/cZKGoeUohXDv6+NZWADsMvYwn
pHKoF6koBL7ERmgFtrwssDv6amiO1ek+MvJzZb+Ua9Y3yCIMRF2cQceBzPcvgA/S
ceDsMLnMex81T5gjmCezU8RFlVBjQdDPfGDQZ+WSRYiRUgmr9EFLinQMf3qc7t18
NFIbQXSfIrBYx/Wzs13skwS21GwY4VRoJd8E05D+XKWg+cLBMPErbO4WmT6dPNCS
2b7e17focVl++6jmz+qgLns4iBuZaR1Eip0mOHlTIJ2/3GdxwAOraCyNPwNnPRsn
vJbyoQB01dYdkZsOp3uKbB+lI43bfjX0yCQM8pgw42kHUHo2BtNL8QlFMSg4tQot
0LwmkVAndPA9zpZODOxdBRoCUM+QvV7N0eNnK2/LzaoWULNSOY8+ggVbnx1YnxLJ
rz6ypDsWRGG1IGdTx7a19aNCtayu4n+5EGQb29LHtdnPHBpl4y2NxRZGd/3C96Du
/7MeoGn2W/OMHVGtE6viuqBOd9IUtTzT/Htp3fffKlRiAnuPwq9BWhinAqIVFXa2
xICvi8fIJgXP8uCl4TPqok+WIj4zZSMaterCwiRhvD37rBapjDPS9+Er8BDnyRI4
QyoiaWqL5VvLKLx9qrW7Sqo/wR98qZxs/yyeze+npJorxSkGSAsjhNifpaom+C88
0xIeihH/xq3f8cxU4RXLi00SUhxWP+3vAOhKEFf1uJOkRa91jUJWyqVUz4fqoNsc
PJok8Z2yrP8ScELR4EJtcrauBiXuTPjOd10HwZBJYayYhffV4GenVdMG2m43SGrV
vSA0IxzMt5F91CueVyG/4uKVc4Yhe8RR3IWj8qbgXHn49zsqyAA2wxRQSCN6R3YM
JiCPQ8q5Q7HHkWd8lRIErca01FnaIL8hzHRWMo4CUstQTyJBTJFIziH8RghVo/Vv
TFuSglf97fRykOd15W7eFgaEhmRuRQED0Jkm7ujyRMZ/h5/up2mEWzq+Nk3U8Pqc
QlIx6Yo3FBONFCyTHCqMgqzB2y39UU22LFfXYrYFiyrc3qddkH/mP3gSPjPcXzUw
2a3e/vm+ItwswC7AkwjRXowJZDWiTf/f2bD8hcprEdwNbHzcKFQjviRZiinMjJYN
U80+Z/6p5/YZvTTGP0D9MQy/wcmmQcC7Yn6lcFvhP1TKJhIWlrKP9PmJvo49cQoy
7TS9E6iNNQ952KoYatGBVVRdJk9xb/LBHUuXwjeEAJ6WXxvxKXaThEJneytkJ12E
TJDt0Rt2EHHW+8Qm1rftj37BAf6Lw2xblOvatI1SmN+hnDbEReZAM8Nk7h1Y5FDq
OGf1v3+1lyfxXRdcipqBsdcf8Q+gI6Y33Qts5OFopuTZBbs5T+682dhAXSIE4TmK
6VhL3bV/c7sZHO3wH/OO+DJ5OFFC6YhsLOpzPapRaQXORXg4p212DwOaBwhs170u
euiKb+6WdEgkuQERwawt9aG5EQsILpe0foJyupO6E2jPeS5rpaI5x23el/x4rDxh
M5rljwT+VfKZN5Qbr5sheOtqeAuBTDvmIE9bakP0UUNlo+KiMqIQtFbNgooDC6RY
Ox4nWq9G5woY8Mpk+on/sZSOOO9/JUiA1kEXg/VDfTIFTXVSzJppqZIOS1ppCXfF
zfQw0T9aC+mTsJdq12JtUCeFNNrUhrSYHy0Go1OVdk213udN/j5dTb8M5XYhx8xY
uaRJGMuOPfKML4+ciUKNfr0OPcxugm4V0BNwmVgU4AnsZmsalM2+GfKKtOT1gPvC
qenwhnxHIA7NQfUBtJl2Dh/RnUZSDTaEZawNnpPu5QdIXrYNC6frDw7dfTOOarA6
dSWDYBATMb97+dfCfII2cQ5tQX4OA8x9+e7vKLTMExccVrxbsKMBwlHYhyzdYdDP
sTZ/aVCSfIdBjM6bGyMkkoCfoWExrtqpCvpjSVbO2kiX4WrJOFm16NiE0C6N2Q+U
VMatsWEasUCnGR6ujHX5fLxMr+jzQi2snr+5k/fRHNvyX1TuXZl2mgc0ddLPEoGI
KKiqLoLzW9pxPXSVnFRUbN+YoaGEZzENjTJ7js6CmHRVGaglLJTJ4fms11DToQes
p+F0mQuF/cXWUqdmNJKfi4ztWLwu9MTFw4AOmkG3yN0r4+ZyMIQdHx+sY0ufmHyU
XPhl3TpUoS23LaRF/t3z/NDBHq7JZtOxdpU8Cd9AIkHxJ1dha3MglO3ZTBliYTUK
vqZmwZ9XKaBu9hjZmKIWLqtbyp3vwjC20w1VIU+AvWfj/HHEMujISRmocBdBpqfF
cq8Kd59sucG44xz4Tktyn+EmwiX4MHOA6dmmpvc8Zpr0TICo5mFGL+awZ3OhDd8Y
46co5WrHo2hBK5hnj8xH36P43Bi+kgyxWYRB5gtt4p1Jvve1po/SA868MdapJA1O
ZocWLX4FReV1pbSfbSGqXsttQa7VoF/8oGIplV8IkmuepdyLFgxfaWjGo0KllMgr
C/pfZI+90Z39BOHdxpWfIzHtjMw71tTZ9sTKjEsdC5fdrCNQ0x4obydaFswrI/o3
7t/ihwgLnYC3Tq35V6GY6o+phq67egeeV4mqtLgHrBQ0Wnd7Bj05fRsqIcoG26dm
hJOpgDapwxowaICy0MbaChaVLQUxfdKYfpWVdfeyG92RPpiGkOpQxcU67pHB19qt
j/e6gz3i0GMaIYgq+nD6TWSVcn9rYGIjRJeix7N46u5/HCymA6deNTG0dVawWL7g
86Mqc9UJsB8MabQRybDRAk7teh0WNPLhoTbARTyb6Xw1LdiSOFrqluGCE2eEh3e8
elTtS4LI6TyNj9nCESFiVCA+W17TTzAiq3ucwfYmcq4APVwbVUDTM7EKQexqTTtk
EVCE7o99Rrtf8AoXYGmkoZbP4pemJtEpZV0EubQiGqbyPW1KNQwv4jwgh9kJfztQ
7H+F7IopPqGhdFa1iiGDs40J1y1vLnE34R+C6iEuGyy0thDnxS2f/dd5IofQAzTQ
UziV4OOFld6oZPv3gm6EWiYLbm8iY4HQJd+C1b5PIqk+N+EMKWP1b2hPwzDCCZrL
fs5AgYpQqtzmr1bAPvLXfdFNBwsRCwxPb5XV0o07oX35DLrfU05e/UM4deFTn3LX
ASkuEl2LchNqSH1c2u8MXnnDkZidTFaOH99hBKIF5YjzJ2quS9ybom1hkOAA/XpC
av1PwMatsgI5ZmF79a6Tu0gzY1M2EvyE+BDGzm3gSE4Cr5k1mtTGDhXzfvWQYLlN
ltNHs5SpiCwgvV6WVW1BbtvyoH5jsoGUbqJd2ILExr6IIJWRRkwazFOdBaaDROV6
Hl14ssk61WyurMDyoFM7I7ynyqFEog9RIlv1BB/sppv3pFw8+EeYanr1pxRD2UL3
Ac3RZr8/0ZmMLwYLPxsC855EXvp1GXtelf1YYBeyns7VMhZ5lD9n1IVdrmQgUAqR
mRdmfNwGaHtlUOC75FWg5GBiC3s+tm2Ea1xktHmaewdMdid3utsLah38vuj7sxLY
maCD/nY27Q1QNqKsuhmcBeXuTdBp0ND8GPouEEqVz0GkfT/un7FQ/ffcvr6lDcwF
Ep6ws+DoyK33tLdag4Yl81srTSg347MGd32/qlT6zWR3u4L2n6fL5Up08+LSFL7f
73zXcA1EOTYJ4n/DUuEsxngIIpgEmxS3sZ/NPkbReH4NavfIAw2Dnmz1BYb0EnTS
CwJc8HHxc7z7nNawEXKCR7K8wQ1Ld4wy4RqU0eJFO6b2dygYzQWj/IHSfLIjloMF
nsi64Qtoqk0E5yoNb9UrTA1gpu5+uazytHVmJxIQCb8DBcEJoFio543wPAXYf37L
SugxcIG4z6Mz35LtOWI0qkbXrgoFRJeUB0KHs9+z4JDNX3Q0jTtwuqqZNKD6ULhy
iXy4dqA0wBisFW0G/vin63ZX0+wtejashppz2NI0sTncAFhDDjXr2ezb/CKfhVW2
+NUAmUiLZ1AccmSf+y1GcCkCaBm5HJUPlOh0T32PHOavbHTEPlzDL5IRu4qJvBzN
plqtpIjpWZrAdRnzzsK76Ytw6VuA9Oc6/rQTSrR9Qo0c9T5OuOjByz417zdHzwJ/
2VDu10GiL+A7o5uPH53NbqzI2o9s9zQ1sUpwZqgJ9mgeRMAFIhGdyWqPKfb4dufK
BWesYf6uIL+91BDhl8xL3fR8uuK5HM4eKW0jpuky1OGM3KMEDDVeAER+QpgKK6YK
rY9IaR9u7IJ9OBIPtqdqxuYMdrP8UvTAaxE42SXfCtuQt74/t26uxFHOzV7xfu6M
wcLEdkssplbKu8lHES4RtOEx5WHbVvJuZQPTAD3WdllNfOMKUIud4Ua3P9w5kH3X
xcgtxwI1X+zYc4KOWNtZ72/umQFb+R6nNpu7zyR6C+ODIzYqziS22COrlN4FeS5T
UkFnT9cG3MjDBGc1TS0utH6Cv/JK9FWTFPuZFfX2hDR51Xa9v9RdKbkecP5PLcl+
IdigwkY2WFTiPSMsQT/0mFIbjfUvhglBilECN4o1KJvYgtHE9VzQ+jCa9DV/wwja
lBrLUUfhJDUl55lTMLI5j5BUd3ipqB0yJ2mJjYpxnjWAfgvXyCuY36uOkTz1lOS+
ansJ5FcAFEOZnFROnfcm9eOLgR+A1Uj6lUz9yx/DBQSuHU7le6MHc2BI3HOZV2N4
CwGUhPdtlwYPgoWla8rNFRz4W4nEVKdFYvWjBQLLnoythHRfzfS84wZrwSa31XRP
bG0DMhlWOY9/Eo/ltOl4+LZApMY/o92zUiivzHLdEtsHmEIwkC/HnkhuCJhQCVqh
sG0APAkoAoClyFCP//f3Acw0oxgRf0/sdHT15hj8RyGHiZyNrZGEPq1+X1RFAcZD
XSKNgvuYcEVaKuldW7OWRF7AWMyGyqogZXkmVhxGnNy41CIOTlI8wOyHvTPAeML2
E8YbQMKJ7VCoqPp7WMkTEeJ0XBZ0YEQIyR02+Wu+sn74SNXV6a1vU5qihpLB1Rl0
6m3QgYruuJwJuFS9x6gDDwEbJKuPxSdnLAIgXpAouAzYir8SWoFmEG22riVyHOQP
Byv1lVC/BwHYp+DmSAkqUWAe7yho8HGfUz2WjNUdzp5IVapCecvBhE6LrPG89jqK
At2nCzi7T6eWDHUDccUZuekcS2nfHSKG/1dxGV0G8lNfpDBB3MGZXLjZ2GV9Br7N
ZoHUvFyhJAip+oI1LhDIp4U1S5nj9sbre/TXOYCj+vHRc2tWJIt22KAde4X9PRu9
c65ciRnor9wCYFkLdgY61OZZj44gHwpJJZnXuWJSfuhaSc0PPCQFOpi78LFFjqb2
4T44Jzgd21ePY6MumDxotNHAMOt/s9UaT5KfE90u6fCUTEHs6waVq8FPT2oy67HJ
x4mVmz95IMEYKOvzmQ1wJHNEBjAElJzF4hIPcDMw0ZFVIo9qKSo5xkqHxca3HexF
qug4jPFq4vbKRtdBNp24VYp5ot9VKKq5hkdAxFcMkgX0eQf2PJcowTaVOEh7xkPf
2K5g9N4x0HL8ELV2eSX0XQCm+NMvGM3S1KeWGvnLMYaNV8J6YzO0igaFgd0ofsgr
vXMP4aeS96HhuHfKomeDXR2S2roG3cV9slCWnH+yqcfI6bbgt36Y5en/OYGKogb0
JsZPQQFcA6bjLmwTt0oEFgok20ZvaLQqsZ0HDMjpZ5NqVQ0QkBfB+TqrZ1TLY+Xf
WddlvAGhwy0cNBjq5MjbkRUtyyIeUncb2j8XYpGN3phqpdP42fUiL1qI3dCaEyhJ
TRQTHpsp+yE8zzw1ipD/V6vOpLMbh6/wVNOBBoNKRkJzh63nMdK+4nxVj+aK3rpM
89EmVFloY+RX1bavA9rR7slznI469UsE7O0TBGP9xUy+HHidfB/GaVVdPS2Xblb7
vNMhUhc8yADwV3P9txbaP4WJRAa1gI1IHnNm5kOePkvVItikGBxzG2TuK8u+/n2s
fT2n5B+hVbIvYxvOB0poDR9+BDqp1xtyCHmMW8BxmD5Lul+H0lmddiyMy7cP+ABe
tRkjZyKeZn88RDF283v9vUma86ISIsDE23fBFv6FyzmN4cdwrUVo5dQWKbhFvsFy
uHslo1s4ixscr8LUSsT6u2ovu8E0t4c5a/lITLR8bSQ9WoXISfMJBECUU9j1AzKm
C8z6FW1v+TAjKvsm/bJ+sJgm6PPDWvqFgMubSuUmZS6w5C6cUDctrkFwrGhCzd/U
sKW0fcWyJVX/E+I1FNPzI6OCj9/frvdcx18AJkI/c0mxXbp3qtudw3okU+Irix48
E6vHkLJyvb8te+tyLcuQCl0Sl/E62sMeX2tPjUoJG2YDt1+8qMBbkmrIJnJbQVXy
UEDb9KDoOv/FNBRxBb1IBadc+52sUu/Z3E+eVNrHSnkFhHEsj5B3/UfVHqEbiOtO
S43ZZDpq+j+DZXtjsD8xQp2Z4c8jmaApyuSeIPiDa7LrmKO23ePxH25eUZlyHtTv
0u7SMzawwHP1g4pBnsqLAisdIJRtQMO4nCijPuskOW+5Epi5thXC+VWc75RvPARx
QQl/s8XVvtNiYOp+e4Anu/MBi+UVszu4/a58+DolClIhdAOqS+oap0Yh9slMknNI
VqBL+Ox8QwtKXyihhSDQWXkpmy4g8Iz3b65P11qhbEF/kLVNmcG/ZkKVqeSEFsNq
drdorAPejGQXjGKN4gR7GffsVhGIw7Ze+KuXEQwP20FYq44b2vy/5iDEJ0523dwo
xZ+QiZ2L5iUpwiSzzFrOmDMQyGTiId73Crofi9P6dqT6qDL0wd3X6aEKBtT4Zub2
BIzg4VNaXujMLG2MnKuzwipYCzO83Ay//jH7XZPA6Ybdh1OEwckKNx7dmWRhBwYF
No3sBYUvX6jos9N9MOc6zvrCisdk2Yf1yvKYHLZ2cbKDIImUhzmjLFdequVX2ShB
DkwX3KCQfMRjTA0FqdyNff1lytV3/+BG8L+9nEOs/JXohwglQWJOIPOlwdJ1AD+v
HpvDwIgYsZFi3dfv+M+ayyeDpjIIFV8sqEboHC18OSNMTcejrpMuRWwjR7NwqFFx
FX12nU9Uj8notr5kqxmGYJi1vdT0fpZmRImHtjI10bIp+R/6U/3pbNLRdHDLGeiB
hdo48UJmZwG60zl5WQ64WUIOv3dyiijzwfyo4CbnRoXIksUwIER9M7WrVGudBntv
Cg8qrJbj5DckgkoWv1/Jt+qauXWcq8KREU6/kMv/iUW1nxNlAB7WSY26Q/LmKwJ6
/7jGgwGvYpD2B5v1jplRea0DlBqrHm6pALwGqyiHFi/120c/Azp0nW7lGykYMRsQ
EOpgy5VoF+GCvrxSuZp5ioVWaDccWX8oX8tV31Vm36q42KIEqKzLX8ArTs6cWG7g
fDqkMt+ys4RiEgMuOwq2oOgYC8LmI2ogRkJ5J74ETXlHCUhwkq+CRZ3JanQB21xD
Yimr4RJ9GLyq2Hp7KBTZAKB1ec39XNeznhjBlPX/KsG1Cz98aOLxDEMb1IBL7caq
a6UD+E825ToQqVn88tp5rBe+K8vtSl1cVIpF2HMm5o3AwUjaO+NsJt+P6wB4Iqea
ZVeA1l84ojLAAzVSsvwOaovlKAY4eFS6D8rb9iOxairL0m6ryO92O4kS5O8hb8Db
uvKKKF1o3X4rhawwAku6LpGRMIZMm8N0ZUzXCwwii/VReulyBUmlL6fPhf3wrpnW
NmS+D6ZWIGjspghMmkmgO2G8VyjP7jPDwuV/AV0QJZeJw5CvAjUAIeCfT7azFNmV
L9zZA7IPDfIhNNxq4NHFBE01oeyzuW8mYqV0NYCZ7qG6FYqeg8JqWTHqXXnI/6WR
nUE6wWoTdBeCEysjxYbjpSWPKgcg6RZRrLYn+eJrUlRQE7IgLf78PVtGkCCNXrZ8
9TRZ1op7cslH9aoBOs/nF8E0JuWoQr6emHDIpMeHfItZuQPIiOTjmDUYWkLTzeO2
cn1dT06SGz5oYSzq7CjBuJJ1mAsmoVuVG+SpRgJbo8KjUSrmFzEs+mnJe6CWMIhC
FnmIzcerQiYXxPDCjFDtci6rdQZKfruHr0Ha1gYXAiH/Zmt9rHgQa3TEJLHuOFXq
Ma0k/lIH20PRnGCLi4+CCnnl/K/d7l3PG2Loj+/fx4aVx6PQQaJkAY5211edzaHR
0Y6tlE/Vxy9/HL86f37US9O0Kk7bRbKtTZYitZAKqhwDAyCfJHx44ynIRCi23zZ1
tIaSHCv89kkbLhN+qWCjvMs7X5HbObmiB3OWFIAxGou6VX+1JWnn+AEQ2HKN4grd
xd9Dqkye2v//bjMRW7VOgCpO7uCwE/QrKoJKgpiqp6ernKUuBgTFFW0Lk0INf37c
BVegH6dBLLVoNHuG69Hg2kXRZ8siKBKgXhYvLf6biXcUvX9oyrcfr4gqSrLyhkPZ
3JYIjduWmu81JYcQyJ1glLRfuUiyR5rrIDpQZcwX658fVE0/j2dfNxA4WvOKsSAq
q/nlSk4rAm3J4Tq2EOIWn5H9yO0zioOCmXis5V6rnPkTEGQ6n0li50K63PQgHGh7
W1fuIKK9ga4NR8Js1DWpdvdDzuBc9vuRpBBRcn5sG2AN65287OL76na4x3QtmMLb
6vTLwQxhkPgUrCVXel4IYmehwBgiEXNzqszrsktZ8w84mMQ2GYVjTYrTCmpfXPAH
yT++SXxl8NB66KojGLn9TVixjnR55kDV4Aojp6U2vKZqcwxsNP58mY7hT9Jfgrpi
H1PXrWgYwjq9CclAwysulWMuCv9Fu1DxNNmGnLOBkPZSIERgzRQ/SIlGOJPKxXVi
7VjfncF1P5RFsCmbp0fvj8hrC3WwDYSkdA9pDMnkppNVEaVD1XsmBic7v5BFYdgJ
zh4CZgk9ZCgFM8Koj9vuQJpbJ1u5vLf+yrH6os9wX21JpQ9i/46X6ZCtScCsyLPC
kUupd612M0ShROyGGTTdODnLFVtL5+cVAq4eQQg6z6w2+NiWgL9+2ZSVsMguPecf
BUpkHP0zyQRr4/X59/OF2RfkLSbGD+TEx0qmS0N3/2AxKpCcWQH2cBKYn+Wg92rO
9tc5thW4NHzT6efDdRJC/+G6H3r4ZCZNgqhGEhknpL5MVPUEgz0APAlskmzDUcHU
lrxCXEAeZnAm3Ww6CgMGsn67zOnz5g1Z4Q6gz4IAN+cILIQKLr9LcabSC8WUKqtN
tpG4o5tmtnW+UeY2lge6yXgmC9PmrKLbk1qyQlPyyXzX5HsP/bDZdUcGkBpHFECo
UbuujqWgEnoTyitWRfkgCaCFxtR77W1Mp+JuwGf4/ItCRsK67Os00eg1Uc5GfSus
0sBee4rXtaUbyAl0W1iPZUuolNwzhs8fl1/hO7s8cF6RciHgjeLM9yp2e/VWEqnO
qjDYy90yyR+IAzAsqneaHwIPgT2pxhlhmq5stMWQ+RkOgTlNJBWOgrgHU0h4vriU
qUjYBX6mqIX6eENW8LFyYaRRTApcg6+5h9bPN1O0JcM/SH0wQXOVnuQ1G60AjW0o
WJRsHZNu757U1Idw60UoB5lPMINm/11annjy+Nnf9LXoxzFwi+bTI1xEstwvuffH
0cp4hBWEGxZsXMnb2QQafscJ7l5svYj4U83vfzbKokADxks4RiNZiRP6bR+4WB7P
xBLMdZfLqwLFv20o+eiSJnm95+BOW/OznNBHtovvtCY0HZEH+ThxQHHf6E4Nax4E
QDWkKgSCrWwRQ0j90hCVXqkL5OQ/fWdJwpkxrP6PII+cOYDfjn9rFb3YLrBmzSIP
HSEtobfIgeaoq8auFTXz0i4kujBWBfYMiErHJWEkQg6DNn7GQz9YzsFXiyn38BUR
LHAR9yuBgawje/EmRo9S9SqleyUdaW/E1b+BouTy9FCuPb/qL/reQ2l0X8G0aq46
XGTwe3iXyRVCvgpJKdIoFrQi838LvuIOOj6Z7QKR79ADbW24oU+zNpKnRR4oemTf
N5lcXp/Sf90PPveDeMrMWgdxFTzdj97I/wUgQeNY8cPUsTUjASn3hILgicJtL4SA
dHzzp6Q3VtMgWIQNO/rrvyoOfv2ETCVYTdZ+ZfjwOBguI8pFTTk7bgXUKdUJyhlR
ugQDIqHLOrJtNd5WznjLKvvPA09MMQyYbIkJ+BOVtqxYWmVMAjIs47VOEYn02v/S
2Lw2i5m2r54FAobunqtjer9mBL+S5EANat/fvNFONWvWW7YHCKTmqGQP5und9zQI
S4AdYr94RwmgGosWqo7vvUhp4ihQeUbyeHGInXLTGrwr7zPsR3+bPNmx7sCH88rh
KRIzYHrxvVq+B33bkO6RiCdsFd0G4RZzzbml4fneyvJ2pZZ5J5oMqP6ZDyC0o6Ny
vkBBmvFi8M8z2jip+hUxqSUrWB3emzRehHCbW4qBFvq358CzC4SwIONyJmagn1LF
LbZSvGUiDqYiZ+Zw1UuYe86vFflQlVBNNvRC4LNHjFHjazAdCNrw1+B4mNJN34yf
JLbLcrELQvBPenREA5Yx1B0JGSQAICJwtPhdOhqrn8bf8UxPqHdmPvQVK0Njq5sg
KhJpdy4QoTytvIB/w0iy4a+EISsK3atLZzw/RXPuQFls5YityKBXlN1zokLs4RQQ
bBIXCqrKjPNoqFkpBZBs+hhTR59UQo8Tbag8T0Rjl7AXYxeMkZtLR2N62ybqAlwn
IXzJKdXHSQnGJNdT+91MSSOaT23RjC7exX/FkuY2a3O9EKuY3XpSpZh5STy8cdj5
e+6QDxQtQEuTKWwOyB/9yjcNKLHUVUIuVcONmX9AmTC42yXUNf97e8xPYc1tMpqS
zxTI4MqLkvaPoRBmKVGkbHk6CSu55zit9nuu/bePeNPyvPZ65K3+ddBSTqpGessh
G12aqtHr5um3yev33FxQsZ3guJZW7JZ+xClQuw8X+iPx4QjNttZoJW8hktL4qLkC
U/H1y3Cnya0AD/8+pRDhXJ7mMcnemsRDx2WTT2ihvgOCccZ8D6kdfTMqBeExdB4d
V22Bs07RkuYhzA3hTQb609q0xriJE+SrpHs44a+fMtJN0tOfvfI5y5e3L3h/7XRY
RhRhL+qNTYaY0RAjsB70jA+jzfWZRUVxKE3LDXLSG1EGvN2sWRFFhxNPTbIlaiZQ
7rlrx5FuZECBOQcbIf9sjNF0YIiVLU8oZLWgf3aaKCuUGJ9CPUYOpV4Thq3KW3fL
FTokp0vIYbezVB7QZWEpO6nGLkULBpYyYajyB3xm6Pl47JfIt8haUpm0C2PcZiPe
zy/y97XGdQza4n4HU9lrgUCNQ9jRY/ygeiPvSSCuugv35E3Om4jxnWrvv/Vk99DP
5Hsi500Ar3Txdc2FIDf0Qah44aMYCO8T3nAqbM90RPkR5ZEqY1QTPiw/2uUCBd58
1LwhoB3Y5i29mYBtCu9NsQDbbwkenHe0LQMmsi0UN8TVQCcagoivtSNr36IVr2CE
1/K7Y6ifSVCSS7RflhVohAK3BTV/7KndG6wq//OzAiq5HiVpGSXs+AfKFPmJPITK
Hn1Oy7LN+xWRxFxwm4dtozQZWCWbqa5PBEHFIE5KI8JA8N+3uLc4FtbqywHgh8Ej
GnCj7IdWI4BYtBee7JMrChJqG9Bfv1SMdt/c0zHOEORXXJCA9O8rcOLslr4Pqji3
cNjcNHnYBwXsSYF0mvQzbIigFrjlDfPhY7RUDwN+HrmqyoXgv9nVpj3UAtMGhzkf
H56aV6r+DhzXCqBiA/O2eQuDdpLF0i0COZpDhxKJBnjnlflIy2LefkC3Xoq/1Tjd
RH5K1RQ+AOzaqIfp9R7oT/pj2AJLq5DI9wqcBddgtTdXZJtEk6eonsNmNVjC78Ub
d19rrOANJ8FEpEsJdTr/JCmvjBBGGqv1OtemU4voGOG4elOq125qsWvUp07/P2iL
8fEUAz61wbeqMfkE2+axGMKaVY4hyQwXkqbJ89yZ8S7kuZguz2mhJd4BlmkvJiuD
bWSQr/Y2zwndVQnz+0o6m2IVVYMmvaWkKBabzwKL3CEPvkUmLTMbC0COZRchHhIv
mwRkcZJwbwG1LUvGLM8/Ch0O3GMwyZMiU39XBzSoeHC0MG4mLb5E49ovnSB5CC8a
eD5rq+zypfcOKsDrzp8Hl3Hz8lVlCTzAveEncrROPv3NHGBEHrKy4mRVf4SLGC39
DFZixSGPM40Gb9LaS5smwAFdK7F+xI93lsR6Do83lAHK7Kk4Ib43MSeAIvXNNhSQ
Dqa0ssG8WA+QkXliX6PGNm+No3DKOfBhpRFjkRTtzmNoEcOGOrwHurMot+WSPmwj
ZO8bF2IVPd6yYhN/CccLOwCrMKI9lQEnENTWt9GEuEKm2g7ZgSBC0yJczSrlXrRI
/xz8RCmc9pnknlCZstrNfH8d9jB1NGk3p1gavWs4NxGsMACb29ZqUoozUdb0YNJ1
v1BbnvnfcY9iqiMSyfUY2aMJIjeGr8UK7a1QE4xX2bDnpisUlOgeJ1wA8cr7mxR+
eJ1f2Q4OorxDiIvjTX4TzvOgXlk0JBkwxXxY0NuD1Tjlis13IcSe0vCCnuuqW0yG
+/PjSf66PNS+6nr6fZnwa7+XsliX46KuhHR6S+e8OYVyB2RqxsGN2Y8do3DREgo3
Kta6b6mlilIWDpiXLbV8ZpD7Qet/Wk3T328GONVbgOfSumDr4k4UjMH+vUbc5c+z
yA+DswdEt88JAtLSVa6cVbDf/1Di0+gi6UQheth5OipsAbH7hVT5TgtGPK2MF4M0
WkhqMxqMdzXK0FYquw78y8IRrXTBNBEW0LYrIBypZlf/CS/aXGLvZdR0jE23lZwo
B2aogWMgHnJsvq+Gd25d197CuSP3ehRp6CVcXEx2iMgMpnSjTA2i5WfdfU0s7zdT
erkqpgE2yuhiNoCm96OWO+kd18hterKu9KCSAqSyv685M75/R18NCIhv7vINVmd2
8vhvqY92tHfSptHejVvBHNbjVAPHgaVV4/kr99ZwZxzFXT/ZjSMDpJ836/Zmu3W4
jXNIS5mkihnxEqnvEx/5b4sgzFlJyIRWsxaJpvUkpBS92Ljp/v2KuVQRORx4Zzf4
8BJFJCTHX5kaEpYm1ryzlDTW7I3/cGuRNVbNue2Ymy49DaU9KhSaj6dD3BkN31q5
RY4GWNS2S8aA5pJuzWqYeRr5o24lY9bN3euekU2TctkNa+NALKmQ+pUXf/26iDDU
82GsQtRVzsGJtgKgXg+Zf1AERcAJnUzKEmsQd+UH0hEUv2DBVvssnAJEpcxUcfzF
plUo+UrHqwpXQVw2WxK2pvs/kbIjvE7QyBz6VsN4fMK+ZmEvZTZVKH9DBl0gxmV4
zFVDVKlO3vjcK18YeYp6qC8CIVWiE8rDmmml95em3elrgd+b0PKyeT95AI11iypM
O7hBlm+8GKyC3WTB9h70HoT/UsPuquNnzsDDSbBTkKt6/8vAUJlzm7TZAaaEV+9X
+5V4v7zDmbDFLOlmQ7QClmNel+m5+edjy4zJWySqLcpXCbe5BzD/fmoOhWHOLwIk
nheBAar27TtfIgmy9CSGAYy086KtkTHVckgfmrBjdyHZkxr/GmZ0ARfScqZjI+6u
sNiTnZxU1wiilSPoN20pM1cFm6t6E9yd10ORnCIX0MdWxBi9biD+t9ZsK9Dc8IgA
NYpQ33pJl30lh4qApoXq00caknobnJZMeHT6N7AzKLtcEG6n5jDy7O1A2KCZF7+B
NOSfakAEnxsKNpy7Vrd7HAn1C3lbhd6KrDmoVrcqA8/4eGVPJ7G90vmO2RZjbQ33
ECltF/tkbVo0/bmOalqG5m0elVTMu0kR1fvv/jCANaMjUfJLSV0w3bNR7+MGAXfj
ycRHQoQqgoOhRl0mLCEtd/Ht+WfFZs+WALhMoPyhzQsAob9BOBrbJAFDZPXHOUY2
li9KopObwU9iYrgCU0MjXUZZLn2boWa/yC0nPA/Bw4/1sNtzEMZHeoFDenm3I08X
4ZArk7nA2hGEMWzV/KrhmUUMCqhuq4sGfsz2imTeaVMJwhraspXSt4PekVyxokWT
KXXXwfYiQTFUh6RoliPsqPKyUeCVOPfqhMQLu2TMz/3Ut8381KbIDlkNz9eMuJr4
esCQPRPXVKFvNn2/UCPFmjgZEEDn8p2H/GOSbIF96ydEgU0xLDQAQIH6oJJKFBuP
QBWBMbLSX4YZp6rrYdkh7qHh0vkvj9hCMSVZpzzNj1DY5KgQBxz7pyLIJwW3DHl6
HYtz/4HsDaPXN+sMsa1E1GnZwrkRxSf2l2Vslq+HWhydT1L7+S3SVXZFnLjhxihF
gMe6lxWNx3mndUETnfUpiPAthr9PeCIgomFYYSEEQWsNWwd2G8C+JirLQIP55eVK
W4DN57Wxhyf3/y7l55dcTSET2aGvdG+a3T8l7UTTpbhFAip4IKEw++dnZp52xgIE
42iIGYdvrrW6bZ7/mPEg0+tjX0uqXdJtmX9N0UotD/O4rqIBlDCoKxuTkVgK/2f9
1N5MgA1KMLL8qfTfCDd54qJLrVfKPWxmjONCy7uijeFISmFABMigyFTJGiCU/yBG
BcgwDfw7805kk5A8Gk4q9CK8x3iC62UKHZFHNzdlAgfc5iN+zb2dTpmvhNApQKPt
2OPuRgzlmWuqFwVhRZWpVm2wP2eiGm1QNk3A6oKAiEiqmhxoCd4tOODOmxxJQz8y
v6QQQq97VGd2yrA9Gk1gd1HrxuEElhgl3C1YI8KAajiofGmU3M/ONEg4lqbW/xo/
QpaEe/44BokkcteDdrO//RE/78FOvhydS7GMmsHWCvXikxXvsuMPcEDVDVoB/OBl
eqHLL0a1SJmJZs0ss+rCaGqBkf55kX4dGvNOYxMl5vRBWC7EjMFzbOUt28uxF7JC
Bq61b3R4fJPKKM8Hrz1TNu4QmyTsnDmPAp/FQehwORWwhtbQAxEL/UrMbqD1DqxO
Ya4YYA6bLVgsBnm7HYRnOfUR+/tH8NdBZPljf2ey6W+DY9TPThrG5JkxVyGu/ngP
9ByBPex5V+BqiGag4k+YUIFgr1aWa/GIjZQzJi+f/HqTgHCCzSDps1+k++/RQQTV
3tAWhzSFnNLhoaoLE4+8RfGH52jonegpvqjbQxxcx1u+FELqRGSCsAjg99UvytFN
D2m7M2eatmLcUHYIWqiCwUDDXpLqxZKwdbimg4mVUNXBF/I+35bGOyKMo+IYQw60
nOOElROStNIzSo8DmnQjz3kJAJeCbmaqj6qApFOVRZ639CqQMSVO8sEwZg6Pd+v7
WDCM/Y5RlwwUOBUu0qJBcQV+eUtPw7peAkTspWibCAwPzA1Uu5/hBL1F9M2svkmT
IyAN05yEqYsshn9CIUq5wgLuKr5uuxSoOs4Vb8vjN47WDel/8FvzJSMgVt4mPRC1
ykbdFeHsa4DMW15eF7mq2MJcp9RuFq3MB194wjZU+szVR3yfXJxhW/ELIZLgshVV
YZ73U3iIk3ONgsv96junLni9NKLbaAkoVGLk/Y9xKlaTRw8VKKkmljewxi6H4dqv
uwJETgxzWkanmaT8VBTVVhGVDMeTLl4b51GnMelnL/8NJQVZZhNxz1jVlwXb6Tr4
YSCFm/YeXsjs58pnIGzAQQ4W5sAEsQ187CplNA4yW5m7OA3J4ThavwFREae07SMd
PrtYIungPrwHZgAa9r3B07LRMpj+A1YLcJrmhxiU0NPp5r8J68x8Gz2E4hp3eVSV
jtmdN58WBnX+HaVUB37GASpRJ2e4NLkNTliZ2XHvRDqFNVp8ngZ7f6jdGdLqW0Hi
7XEQ6Otk0J+5zpxpk/0nn24RhASo+dP2wKxrnmFEpSQ2GGO0LKkRNuzvN609LqqL
Jk7hcvJ5UEDo3KZiMMERPE3yNz8VpPG9wnTEbcwlXf/4xeSsjDwxeczcuZDBlUsZ
IG50po5qFgShELPsgmEKw3i7nOkvSvkGcG55ueOzzcmFaaOdDX9YxpcQJbdh4MPD
aCK8yM0LujxeMMzybUG9Py4yvyu6gnshuP/tCyRABcPt5UojtNWqoQZdD9FF6YXy
hqlDj4cs7ng4LA1E2i4ZZdppXGYOf9yM19BpVmVozEKpINeld++hGJesa44gq0qe
sM1kAKeKz7wDoYQ7JsIzd+BpDJs8PnXxD3sXASAi5w4Lef2dqxjwhvi2viWbid9U
u7bkTln0WiRoomxuhwhesC/FAwbd84u46De/KP/tU4Hje1+ICxoaYLwnPhtW2mb7
3sBta34JwISUVECldRftm63pL4/Ic4P9DsBQG95CRuCq/W+xPP1tm0Hkq5/nb9pd
IDtU/ozkT7sQHQj+07D3Y2j1yAOWthxtWRaKiAG7g4vBalrOVBD3rS8ISBA8IW4w
PBoCnaraSVoIfm+r2b/8cEZCwzHSYNcCDEZC1qCJgWTsxL8HLA1B62Q26zPs4Fxl
jEd9tjwXdKU2RmixCHPgj6lJVkCffivApeBStK+FkzxPGWhsuXyWTJlSa0hy7Vpx
H3hTWWs25xKwIK+7k8OqWaIM/HJ3182utYu/Y15/N/px76PTV1lpt7PqZXL9TEbp
bVDNVrNOys85ntdEZe8/wXF3I6zVyp0KqL70JfJIWRRwB84EOpa3gU3hydfDSYBO
QMr/TFx8oXuB073p3OnklvXK0LCLrnp7qEK2gG6im93Y+7+B4SoasjpmX7ROqIi/
mp7N6a5uNGIdxeTqcE1UEylqpZGGPB96iiNii+4C6k0DEKHhjSYKKdt2Vd+cODHA
zOkTNL6EXQ+5mvtg8ih4WVisQCECJzBXs3II3eXtggVTcC/IY+XLJbIcB8NkV4vb
xybyCZQJliHAxQROR+M/kFsqXX9IWkppohufx2d66SmeP2b8kI+jGftCQLwFdoVm
QUJxC8nLGz2FRZDAaD+d1uoyHvlcCJ+5AcRsYudkDZw6EXoBIDghl+izigyeVvrc
FfWXxKSsXhfHFeKb9+ZlgovI6G+0hGl3ppOdObrKxoe5wigAygr8QexsnVxCTCXD
hSdolqzjp49DvHm8tnDBSp2r5KdzCpan7tUn/sM6+U97rGDajC5Ryr63ey/7Gnjm
R0YK1MDhUnTQFhwYmRvWlWeACBR/kVsn4UwjrlKygcq6OR4iRQX5vS4lBDNvc3ZG
Iq1i7SAxiVmek1xvhXBPXU6e/EjJ+4wraqXuFxRzNgQn/HPypK1j5wtZVBFf73hy
FSXbn55f8u/6Dyitv1S4aNwNkCLU5NA/CZ40cLVqtGrsC/XeAn1Bvpkw9HwAg35B
GTX3wjkC+rNSOqc5X3/2T1cFj4XgddQbIks1K1Mje1mZN/QYIzpsKBl9AWYgbsxB
BwkZaO8t99VtG9veEm7mR7qXnBQJUDiBsifo4kD9opuWocpMinLxeaFNzRJEovqJ
ignhW0IT64wfFWEVsJb4qILb+i1sjFX5rtQQFMmfiIjExGKXvg4NAPVGrpHOQoQt
N7yfD7aT/8V0YoCZ+nHAWGPOUEva1wKtluGWeTrsWZXwHXR91NNJKOQYrjMj3ZUm
iErbvleuUszIdauNHL9KWpbaPt77vm7vpiWCKTIWdw9x+elkyiGxDLklqgNWhX3/
5OzizVjGbegkANUOf0cxfoU8n4gFAFPtOLODJU52Fyp0ukYJhtgwFh0yDc30hBMN
vpnPezvwYr2spRsWjZBsDJ358vXMAKijAImGwb3QgFdi71dx3w8vGhCCLVqjcWuI
gerQaAhEUtQ+r/TuT1nauv8I2N7PGDvdR2Gw25ZnRxIy2XGzE3u3HD0sX7bajlAD
4/7V0jy3o4fxxb32bh94UlfV1kS5E/VDhg111uZdLuEWv/5/iAKyVhljOooVC/oM
sdscxHfArqn253kW5mxwE/KIobSOB02uwgPHyf3j71M3MMyyRSq+1qNUS3TDUFw3
QwlKwg1LZMqDqDM4zpNMJ1ErjDzGIB4NXyPKS1U+XcKOS6XS2kPOj03kMtMdFcyR
xmtObT2fcxfnwW03PwM122ioQhu3ESsExKtf2CvHzV+GVqmE5W8sZZk74vWxs7Vc
DRP/E9LMxjcg8lZrJJZAZUXvF2Pr1j2ci+lTKCmNsSrvRip0opC8mJqWaUQH+8aX
0X+O8JD6DDz+Mv6r0hcETgAHkPF9kITGlihULas5sMGfA+Rp7kwIFQhmRFtPR0tp
1f5YQhYPiqk2qSZcx/de7n6CeimSAOt3hW0CXsrO/wr2kX8QmW/yon+QQveeDZS3
UhgUrygkRISRwZBnpnzpCnt4syxG/wr/yhjuQoadO2tLaE1HLp9hJW2z8bl+p0Qn
tO2/wgjTXWbLzGBl6yCd+oVYzU/nClfs2VzdPGIdzS9P23JWM6JvULfeanzfH33T
Yj62Q270Dbt1N2Y3ym0eUuBmfB0TsJBPeh0VnZ2L2RKD/L7nmZ0Tin8kb5aH+v4/
LchaOsFrvZmHrFrJfM8QuaqhTTUMzh/NPQ2y4GSuQxKnaJRrlEoYJai5HfMnH++s
Zt2afWA8ojH+irkCzcPVrQqqkZhf9ojAUY20gLzctpqm2gm6ZHKksreCKI9VYl5s
POiBPDQDrnP9xIvzplbBTkP/nN214Y1qu6r1ycxip0TsjcaaurkuSKCE2DX9gP7T
bxBTYW+/r/ax/KdXav+qu6uI/GSMAGeES6D74ddqy7YCHPlBOoN18sn/2Al4Yqbp
nSJY0UiJFRTuUyF1TT5o+1QjrtDi0MyhhRdcyB4+80+5cOuwmyrtPltNgkB7/GNv
qGnaphlrnTpcJWN/TnWjr+uC2qmSKCT0YePl3WJJTnPteeN2rIXA4hI0k2yBMu0A
YvWIHCfqHJDXL8MzpVMbOU8CsrYD6BfaZrON4TekwbPbS4bp29p2cGjn7M/iTBa5
g3WpftfDb59IPnXN8eexxv3TVPmxU29S8sCHADPvhjO2JUgfGdne1J3qMNdvB7l4
MExyNzktv2odEjjNAPA/n1S4GVMTgz7CkLCkHjElUQy25rSISiKJeCD5MAIWUTyA
DOuJfnLAVVzLtY7gfGvzSHKdvQB53NXga6pGXO/0T0Lhly3z807Uj6Up5PVPPUq4
O278C6SNXqJLlqMHm3i+Y1CWTYGGeOoO2itT7SQA6Lv5ygz4ZeCAio1UI5x2Z1z2
BkDc6BfKwqeshonY3KOAOWFjXi6iG08hcqyiVq6J4HQkpgq1yoYqC3tHRSKm2oR9
MnGmE4sVMIgNpvLf5m3fr6MuJsNAuljHI1i7TaqfhelrLIOisMd0KVv4kCmEMuAI
b8TeddPLi7uO1t80aqOyU3X2EK+fpVyM4MIFFJwo88dh5AzzIe8FcqdnxLv+TYl4
JEIkWdmXTm7n0IuMKoTTpmhp9qSO4xXaBZkSIVOcImhih6/UuiA+yJjcKFUVPHjP
vav5FkFP1H2vNbcfliTL5xQzhFf5bwxDtdPollj01eaXm4ev1+Uid7QFOD6q373u
qsdFmGeilRxH97cy8GGQChiifhcIpULH5qUiDC+/qmMJurIgZWqF6fQlvIR64YJq
JwqH2vzHQ13Q+c4vjXl/2qZHoclpJgDy4JcNGkfcaL8L15Ou5JPDwnnBT9JFCZt/
vssiYWUg2SYPWIM7zYA+MrowWa4pOU177DxtcI3oNAfOazbxK29oSw8kqGMWwV7Q
3oxajDG1ytazsZ3Ej7B1ZvSXXWW9sJgEgn6bkxcX6h0I+yC95/ByVm9W3sv2CP6d
6OJZ3eEQP5pBWqLBwu4JgJnfh2/P6sybGMjr8caTaRABXKlKfcjAiIApmniQ+PaO
ZBkfKB1v+ZCvgZlIGgU6tNJW6xPPlkcnxl302zYYwEDSnXjmvFCq9aNLsXbpKW7U
TM3GQmuTitHI0b0t5oGc1Zlw8L5qI1HvAx0ChJ7YBXjb47Zz8yrLzDxKoqMTUpN2
2wN37WiMQtKk3Z3ei3ASxZwmQ36ft3GvtvPQ85Gl2yd92X0ClOoA1U/F5ACHrZE5
wb4v+HyXOt7P1mj+PUiSlSoPLDaZzh0lzrvlRSISfVIpsYYtycwsP7XpZOFHaode
3nYIoW9uJsa668v5rGsG5gSDoIU5ipBOAoXOfREU5pqajE0tYveT1kjpgFGxc0kO
ZvvJ+rfc9vIiTdUevPFQFq0fBc5h0SHmIro5IxPQ7Tz8LADLN1WgBGDkgRBkPUML
TCRILrV2Mk6G1zCIURnlDHsxh5FzU/OuzOfoN53UH5ZidjVulN/+IPzjvbWt3fho
QQGeDBbRH9ZngJsX/zWcN2X+BZy4DX8RLFCJLAfZSUSKCJ5cBMAsjzlzxN5OIjfg
mHSQJDXKNRSNt4EJhA2ab+4yAI+bYlOrwZQlvGwcLfL1SwE+y8sFFpAuEba40Fmb
fPlV937mDlawzlP4JNaHjFhfaIndIvGk03drKeC8I3VErkk3HrdaE9t5EIhYzT3a
exU9R6/M5TvgyWH0OuXxTrRS0hPCfqsawn5U97K2JfC72H4JZEhMY5g5fUJ4UryO
xuvVO4zS61/nG1HxjlMONNSagMrZ5KlWzdCyb8nedTH6otO73jZnkdIuDw7v0QPM
m83fyIf6IMEkDNRjIOiBztOcB1d5iLx5Ujrrj2XHFQbq9Wac3vrAuCsSJ7oTu3J/
vegJLePFL0zy9k2GeU7SJm65rXoynLTwgo9Jxh2RcvhJcXIUBJ67thjYpYx7S4ON
ViK1+MPUBlZ39GoNds6P4bhrUyrzXuPPKwfgLHrcL3hCygY7S4vahCeArWT4pNeI
g2UI+d9NRm8EWZTXzvy8/1kt2e7j6TemXhIpHhaDI8Fw6QcswgYbH56eH9JqbHQk
fRGqbZzlOR9zOZtx4DyNRi9kQt/tvl4oyEVTXZ/MMaaYyIpU5Gofs3utjnzE/umA
bkUrjxiI+KMzOl9SrzLY+E2ifSpA2T42C96u9aHBNsOQ/LwHGVC2c6b+Kg+SMP2O
99OuByVxOKgZp+uH6AV4KgML6y6iQWR5DfUfCYmOVUfiTkOaREUKmS59MqxhFYip
29A/sE21q/FpTsi5/yjrqWs2XjQcz6N80hjypv7hwtsEGHAOuT7O/lmT1DK6E9nN
jUtuFaH37qFTs/U4rUPF+OtnkP7kwHZj/nTL2csXT+0v64mNH8yXAktBZ1FtN3JB
dY1Idw4Thit8LpxwJaVQxXOyvUNAmMSFK6POc9AiOh+OBOjd+pwDhokdz4DQg04S
a1+f9zYtHBdP1VdL4RoOWdLAnfgx01KcWvsSGqaPuXO0SFNOpdw08BPcNBs+2rVA
Bk28GmGFxaP/mgyuwGkdm4hif8Y3mzqnCx/HGC4SbdmSxl8TIVXopERgNcR4i0WY
tQzZt01RREGD4an4oZLVo6NVMMHCE6HZkqnH6lotYu0p+BO6Uryyw8yMzkuR5Jiz
TEE80HzLgju/hef5SpGgvktWVdzQx+LOrWZ1Hkfzuvhgroq7YE7kqMdKwA17ky3O
+m9LJessCM6XBaKuwlOx1Xo1aq9gjv5AnnVQBQakb0croZkyXlsdbJ+T3u0qhKTq
EMKxpdkTqkG6xzv+4Y0kDMLKmSvArSdKPrbU4adiy9kbV4B/4vE1Prt0K/6GZzKT
54F2Cj+TsixjtZZHF4YtOll95XK1tjhUvYCDLZXfLi52tZc+4GWOFrHynmDSsDZe
Mwg77Svlk+mfnwxo6WeFK+qp5qVhs0Sj4jLuV2ZdcTSfohNZCL3xaZ/tUVTFBCkP
Llpi+zvVwQnkpl40qloELPFevvWtiSR15EmaivQbwfvEi1TfZBRFH/8rvXHtDn3r
tPxUxMO+4as6VvXAYg5H38ioLDvxMc5UrxxBN8/Z2oCSI5bSsdNcPJ8sgq5YYN+R
C7nUI+oNARJgwWjiXPN7T0EXM+hCdoPH6x0UGFHqUL3OK6/vtPutVXAX8Cn57PLs
dpC8Wls5LGASQDCaQWj35jf8Inmk1TWJCN7urW2+4X974clWLtD5ppgH3i9XyzNO
Ti2Kw6f+Kd+7LLTkwj5tryOvaemXep14cY/gPTJkh0dYopUP7qROIa+fIR6rMek4
mrwpqsVDPvRor+auJDTD3aPHeRyDIlM1xM74stF3tss2Q98AKh2qYVoteLhUCaKH
UVpHuPmAKkPYXSHG7ofiaF7NBeIHxVx1+mfs9eFZ9NjPaja9pN5gHvy0OS93hHsC
zgJr91YTd+MBkl+huYDZdw32QBj4LgGumD+rhHiUHOiTeqr4aAGOYZxS8dILV6b4
sZuN3ydIlWypmfZthikkvZFC/Q085okXS3MHWKaMXtbzjH+nmQVsMqt7uxSw7oxV
77pviSd3BzP6gbZ/DKyCDl019vEvBkT1QylPJiiXR4cihvMgnHuAsOHg9Luvo6n+
yVTMLETvDJydLhH9doQCw7IvayG78Ss2qLxY4nFRPeEhX/IVTzeblH6SbstD9BVZ
UYXFubnAM0dpbyOVlgopoFgH2Wjgwal7rSeaMwMsKHCxzrv/lP9hhOIjhSs+diz+
gseeTKTknI+g3AJuih1Tb8FneOXJa6N56GZZyAH4iHXw3Phk3pLwvxmJZSeJ8mX/
YlFu7+XWWVrqt1m4bsW0FCantYqrTVX7IOEhydwS2koUaUwR2vdyGXqloMyX8T8g
HlrTxMuj6VQ7qAqkUw3KHdcBr2NY5eGM0xBYGKq5TascI5yKfu04DrDAHeUqeSaJ
hNqcSpTLcqnCOxuEvi7DViQFSA9r+dNV7DSZyXPPXkjJXLkovsRTz36V5afxBQuC
uWZDIPHhPcHfAoFi7oRtfFU2YCaBa2DVMt4BIDhND7qNPFbDBUY6Zampow86zd4I
EGvsIrwTIUJgpk0h11alZbInFVsXfF5O0zxZc398xQ4d4OAO1yukrWAUFckP6rYO
jyJPO7NW3G0fViSGnPXrQIwB6cK5kitz2fPRah+qFeHJIcROh9f66tqsuWf4cD4h
tU6EJhfxBf9lUwv2Z4qN5KSSZbxGf7xitDbVEY6r6IJfcfe/xHTBhvE6AcIjaXeh
Fd1sjTtBP6BBn4ON39zWv/5KAkOs4VUm2O+xKhwq/jhBGWuz2uQ04ywuSQMqy5jX
AA048KNnIYXHxgIbfK79fBppuRpOCD+SohEbsMKaC13MIiwz96QooRyg9A4XnyZQ
WWOWAt4eaIDOOv8UPuZ/FnMCyIfNbhCkz1OuRCzb6c8NkLw/5A7P44Ljdt05ER7V
QHoPzwsuxgeWzXtMMkWHHRQnztavGNby6m32aBBwNCs9ZHdsreuha89KPiUyl8nC
/S/ziaVneIulxXyFGDGooe2qHFfGH1jHk7rFE2Ed95HOvqOW0BRhIOfdojcyYZQO
dClPhSSw4R0LV5hA1NM+4jA2Lk8uQ13RI7Z5UIvBxllqlYJDlGUYwDWOvogMrjLy
w7CJbsaqWa1TT1BxzGyUxE3VUAflJS7OS3qlkWrDgBc4Td3r7AxvpAfnjHe45mSi
24HmBeBdqTXQr/hMzQFVP64caWB4hBo2UDdPSBSIKb6+B39vaUdVl4UsNbwkhkfS
qUfEXUxBEB7RLH1lZxjVQ/UUvx1HVQpKKp0XXOXdwgKyaqsFOgnZyorWA5PDTyFP
xOtK2wLIgm6tVYEmPqNHvMUtHnna5KH1bFD61FMyiToCN/BmW7qJPQlDHu2IBguP
d8n7Op634FHC3hwFIR4LpXGnefAo6gs6BVA56cGy9lWx1iJEUIDUMTxmO89tFEOz
gSNzeic4OlMpEINC5I/ZATIa4aMIaFKEZgK4CkNwL6Z9zHddPDFWvVskJORYIOap
8hiXMybaO1Y0oVr/fqm90Jw94bSt42UDufTEf3DndfLbswQP1PutU4OQDFeVTm5q
Y146V9EX94CdQhikZ6e0fPhQnVwNB4h28z82wP+MOvBtNLcnmYIJtVt/bB2oBbi+
Sblz03NUcIlara8KeH8Vw138wXGtspS8qbUqLJ+iq31axTHNJJAR/B+3vrlJQ/yQ
fFL3oSB17whvVqqK+0ncf/fe5UAsZtI5QjDkW7LjJCo6iXpUJLxTd+Y72XmPLXLE
BKkUjYzqO6b1v1HAuw81sfRO77UOn9FgT2SGkh95JRvIzN4jU5WNy2IuCbEMVcvk
gAhfnAAbu+WGmEXxqJGMYbArVl6lgpXUtYqVtubXne+5bizIdDQdrNZP37YTx3XH
dCTmhdajtlMqMdNxhV49eOmV8FHCCJx5W10cKEIhllK8o3SeMaSvtcLRUi/gOIOe
IgIXJDB3e99tQbx7FXWLe3dvi/Jvf3MqZgmMVmAJEoE277VKfyw7Tjk+MT2oArAi
Ohuk/cAzU5LvJRDbYd/J1b1uFuNSyKSYEVAXmPvOaJC1XQ3Q2aX55E3uZUhcddry
j65xpsqc30xqaU3iuvY9nNX+yFS9SjBVyz36ou8g650dccpgLijWgm9FkFOyx/S6
9TnsLIO2es82uuWSa9SJF7Uj68OtWVtSHuLJKWHFYaG0g4tDaW2H9UMyrS9X1ivW
duIassr8mEG0NJhu/rOSQhRlUaSyPDHO8NqwRwPPoqYiZlefEP65n1/UvaGAjZIr
64l6LUXL5H55577Q2CERYH5EcmCgN3w79nabt7JeBw4pQGciN28DPHWkmeaNboSh
Atdj05DnbvlXukAY8WilXowdleLrx0urE5XvVnhxt8Zu3vCNmEoz13ch1itfwzmA
xBUllhxetYZMJdTLQoKBddCRF74GyUDSXr6EKtZC1xWi3N9OF/0eI0FrP1q1mdB/
+ZqaMx3YBShbddsTGhxYru5+sAfIpk1ZaQh+G7dHZFxmB9fBGEjS4o0ilOmX/tDy
BmPAA6TrrE8PWwMggbyYX7+2ecflptvdV8IPGCo1b2ul7oI+2fi+tKv3PUNbiyMy
wjvCNRsLQcF91YdQQt6x3bTXpMiaDNsh35BVYHCwUytFAn+Ai/Yq4ceo9L/ZOLDP
su3+CppUsPePBnvxas/zDulLkoEAzyo8IroiHVGE1QOQBqRASRmLC1AD7fLSdVhq
GRgy6Ar3OzOykfYDEKawlHjj7TQVQLHJH/xs+/y+pJG3cIyMdgACUTBAawmkx005
g17tNiQFP4e8+8QGsKwQCCSldc4gSb4yJdQZZMezWnuKuMc/9T19vZHHkz4FIuZ0
3AsxPjMqoO4DJyTYldyOiW4qSUDVlm3tajlEv3g7/6vETRemuxkV9fx4Fge0P9Dw
9evKsay8b5vPtNrOnPjspqGZkLYOo6/IGD3/tEC3ZI5gNsWH6511Q1Gtgh3uE25F
UTUw7fyBTametHnI2qfCQIXjYuP5JHrdjuGPkKotVgRhelCUzkIr6vdAEWg8JYeY
BhscdZ14D5ADMxHbef9wGNen6d05HJJ9RjQeFALGvyar1ACX+jP8JgakXDMYy2+g
9+U6bYPOIn3CTlHKOX6MyBCn0gSPl2GAVcVCVZmSrmCv1OjW1yubUEAvl26qI0Mi
I+1kFh3EpUNcWIx53ANJ/05B5y6bf/H/vrosmYUDBT2oNSH18IxrPW/UAnmwpYkB
o8LPnwCQjP7Algnl2leoCxDcNO+U1RbO2dnUu9RDCzfzJY2WPMb3o0v2UWrhscDW
dAL+E8NcaQVf6EGrPyctuN2P/PTbt/vtaOOGgnpM4NnFxfc1pPm1WQW7+5My9hdw
voB+sCUcQlLs3m/WVjxbsd1MPoXqkJ0uvarKn0WsrrcCtsk2y3HF/681f0OY27J3
GIvhoenmTyqYwKgqf/5NW9ZTfu8SC1RjOgWRID+yEkgLkwwwAUpebtyeRT9y5RJn
p6zXrjzm+qDtkSQxpTfolQSHxtfdE4IqGKT8L+1TkpitKyWDV0y2FhS6EhmrOwc7
+Ui6qeQfW1C5TLl8G1iUn74i4iWqVx0p9taVn/EZb2GYcqhQv+xpK+SoSr+FbAjz
n4orAUa34WV+a6vUtDf8bfX4+nNSe2Be8UT1cyKR2W1ZoOk4i1kRH09MOvZVzICZ
QY6kV1Uz/Fl0nrkQ7IkRCdB650MVV2J31/tZMb2bx81PisE/3HrUy3+d9RVCe85g
XN+218m0rstlK0tw3MYNBPQ+Azu7alJ2AazBafH7B+zWmYelOTvYWpED+HOOKOw0
5Lk9fAOXGCcsrBFWhaOemN5jPKioYd5ezH2+Xj0el5MLKkaeZTeI0b6iryM8/onA
R8Xk25fVmVzCj9IihM4282n0x7Y55SqMAIcGe1LzvbaJBBL4GSuz0Rry+VSS2B2v
zvBRJT5v5sKbxrCcyfjvy+OIOEMtAeeQLsnacOCqWoiqsvm7sFX10a8iS7lLYVQ6
TGHoE8dEptGUwItl2fVJccuGEY8287LM2SUh4G/gNwCNT+TPmoN00wZsoca3H+YQ
mpIq/rlbyyvsYSy6nL5iwqxubG+02d1rkWqr+s3/qy2cys3OhgtDZRPOfR6ScpgI
IT1X59kXiNc1DOLGa0lryuxEy+ZqM+peFa7b6OTDpwtY/eSf94Ucq+NiqysYhfaa
X0VMLNAjcJl42FBdRpjIbgkw395Nmnf8aoKxeZDytLuUwWkprmUeG7OyYoxNKRjt
1iUwnO6L2FDLHbvUc7XLT3AWsYp45ravvuvYoeLRQGgEYuZsFGu7jpseDG00WcPV
v1EMInBb9n1yU3eoOHNQrtYsrkpRQqwYdhNImZBOfEY1vbPC2DOzdWDT2FW2Ofkc
yDSiTFB5rq6G1wWaMFo2AvvP0V0uctFZKI76Mo2AOwXC3gaqpUBUAjZTCkZfh8T5
V6GThF7uHNWkxTAaIOZ0njGuyp2pgomtSAvrWW/qr/8pOAqm05diAKwY3F8EI05h
w4ZrHpYWdzlxMyIg4h0tdcu2zE9Hj/7fnIOD5T+ziV/x+S1oaA+Ub+A888EdViAi
Pwicr+MXe2X+CXAOc3UfukOPTWF0qToLWv4m9g1V6F8pxjc4xNXk8nEBzgCDxbD3
70majBf+xdeLtu7jLicTD+9JOwgzvSroO88nGaf8CnHQA/Ywo1zCyEAcjtADXN3m
AXEGuh9fIqvPqA2WMtw+PNEbzI5opsuzNy1et7wIi+BJghw0J+ivDc2oHlI9X2d7
BhsimymX3/wks9dYqmrDIevLA/1pNEpvXbYvWBCxD94P+xKcXuVxffL6Q+t4d7pj
dYz7tcIAfxJNTaJ4iV9TWQjrtLbkt92h1NyHSlL5v0ZyPcF7kjNiAtUYDgEQy6iS
snrcbYL/07woQWpF+2r+LNLsTCwer29PMguFn3v7oLdfgqG+TKorfYnPJ3Rb8cHG
zRqT/Q2UTKD5bqGn1qQfNQ5JHXgzkzf15Yd+XU0KURhsAMx3OScSSPUfbqENtmCi
dzQZaEDF/ArepEFPECPgtePvXuDzr2fEvVSN5Ffkx0EkMHT1K1stuF3sSGQUJeSx
qGKyb+p/jMrA131kkyE/03zjQmL3B0Y+joc23uzKVCcVOz4SedSm7eTZ7TMDrAli
Ix5cF0CfUNuClljO5ZNq2QHalrzRIh+2mF6z9fG0+Dkdi3hYmh6bLYlCMiUfdVoC
wom+PifyPUWBTyfEfOOH/gsJG3FzHqhWR1iyHHrGJDt4oyNyjkUqyCBUcTpNLjyR
JtbCAvk3VO6AE1Q37Lq8vWvmM5AwKcVp7r4bDX8MfCL8X6ykaTiqgWi3MKAYFQMN
OglRy7O6Dcm3rxBIVRMC/1Uki1T8QuILaDQNlgm5PFek+f6kB4mZ7EMxSfoojKnI
mjLuHDxuoc6FvOYUmqbHkRguo45N6DcwHfTkeKYgJfK7hTXj0hvcCxz/y/A/I2rw
D5mScCrvRjZsV1XKyVA39yf6Mz5ZOx0H5IfNMI+Xe6hmU8KbX5Hcj3BR1KplCz1Q
6YiKf79nH75QhyB3GjyPfxGto2vgHBbx5zMc+YhblY8fT3pnjccnnT7tvbdTreGw
a85PUfL3xGuV0pKAfbj2sp8BdZPja4GWLJ8QJmujHc00nvvjPfsxmz/jT6Jawcbx
nbnMUPBzbsqZAV7dk3f893TrqRbOOQaHnMXe2xma1zYSMSM2OAL3AUmbknYiysJf
WbOONpeyHlfMhvinsT7rsndqbX+OP18mzTPzH5LgVkid+gOhShSDJvKUzoLgKNoy
i07Js6PW+86UK7F2GmyeTd9ucHf4aPxr9sRN03ScrYC/ce99tnQGXe5WQT/9AYQl
D2maeWXRjwi4SfgxqgG/LZp3UAyn1MXCd9WQXHcRS4V3XNzd8fz3XdeoDsEe20Vb
lMx8WkikLR4WrQS3cExpKXkeZd1eXHRrQGNTIdkEHMqpq9P2+00DubBfTm77MYCa
an1xyOkRTB8r9sS5q/qlSUvNbJC1giBZjdhsu8uFAwleLxZZ4CcYr1Ry6mmNbFu3
1kPkGJFtxkSApcrO2odc6wnIzITnszyXxCCPcE8rPDktkzLtP23C53SqiEy3ExkZ
E0sS7YP5kZ0IZD/Rh12Isn7nrtDUdcLcy3Pp6S6mIJcn/pndQ0AFnqzlss3viWQ0
H5bTiHR9x1LfI2QZPJugD4wr4QLSkRHza3k1p0Ps5+bikEag9G/3LMz5lNI5zXT9
aWBRi0gWlcmrON5YzpOepzYudn0a2eiBijUfXznlNqx2SxrDJYj0hR5je8swBDhZ
qv+coDuQXkLiIhE3mRbm+67Hfjw3gKOkWdoG8EsobFoLh1CRkKPJp7HbL2vtNxmt
7acdyMzUGMWIb2l0+LOh8Q5FDsiAk/239jmUcswluKkEqTzyMMx9Uad4S8P7Ux9a
whaeYbm2ObYSFaFzKiOaXKH3DiQqeHbaMUlsmCc4XIe50GLADcJGkMNDAWbDW6yc
BEhql32sHJfvivd45ouNLHZ47eG6NyPawCrn8aawkYUUlimgutC3Mkd0mPgIuEqP
60i/b8fNH13pm5Dr45YYx3y90zr4CVi/IONWT8qsVsBi6OnHjSqRrcC9rZyePaDb
VepA+n0FB+pXkAO+ZxDKGLznGRz62SGKl82wqiDU+yMdr4oM/83QwWfJIfcFdb3c
vICCuq9fDAlD0rkhQEcIMR3+htF0tlAnA71Yb+IG+la7XD26rYREapHX6FJV95zs
AjuScKvnAjBhya9HGLLu5TqQPIzXUAG3sGD0ERfwl7VbR+AStqR8EAhc/kXhh6eq
/YaeYzYuXv28waJ3jQOzujq7zRNIjIIVSfSRyEbbWM/jWZ02HlsNaS9PvMI2cj99
JucNk5mg2PfoncA38Duf2+iO1rENrMiSN+BpJf8WIPe4g6nEa6qZ6l3o4ZJy5eUt
yHOn/0u3r0PFsSXGS1zUucSkWB6NiyiKnlNqRq8OdraYvNjDElPxzRMQHm0RQlMy
d/RFMiujMzjk2YcjzE5nmdxVTFnIJPQrZ8FivjAQtCswgiu4HE6XxXsspqxhrmo+
2BSQ6c6c+GyYUglmiJO8aqeFj6MkmtlWt+HShqtaOi0Y3uSCwFaskXs1HXq3sGqx
NJWT/Eo+Do2V3sTF9BIRPM/pNSrQxz695DmVPmjt+ElW3qAQD5MkGYOMx/mBiiOe
jPbrP74XWDl1xSjoHbdfT9UsAHdwvOlh4yIJ3B8k4TTXOLSZ98d+okYOzKFBq+nH
6iEK6yVfH8INnaMEaQ3y9Qh7Kqpt1yhgRL8o5RBlTCM7Ar151LRU5AgYsrS2UkAE
sE5//xFTD0ERlDH4+2pTk69qDwYBC2Ri8a3hh2NNmP54uEOcQPCw0PRn00uObEdl
J1eCXg07eBA4X5uJrPd6oNN9odLhaCF/LMuvTUxS8Qo4RUJAi+j9ShCPZ2CN2L4/
WHeohFZNttySmxjuSX/u2fMUrc3rGOfX/hAWNvCtOivbHpeehF8c4bzl7TROHdgc
oSTKUeiEa8swcyBJUwozqh3zL+1Npf74J6j+44BCX6R4psqUYC1arT5OHQvzDlTn
69HH5ZMTVKbl9JWUhweLJGQCgpGB1D70QoKX+MwzxeVtK2zIRCizhE0nJavNtJm2
UDCwhyFf+a+ZEd+kiUUsM752PbibpfsiVZQYxUnAibQnBXZifBxsWf6FqonhUHGu
FnLZxxvhb7GyGUG6dBgQGBBnFqIwJk8w7kmrLbxylyizplGUpujhHLoEb2mGxJyF
RsEzXp9MRrKmZ/uo0WT+DVAET++JeV2szUaJZiVPDEGnBRg7TlK1CHyJvHYZ3WLj
9CsPknSdnksgkCpRMCk8p5PrA9b99VX/UuVqkJ+PX+hxdHlQ9Hll+YZXi5+44eCi
4/UpL5R2deWOLUcJqylJreqOUxRxlOKNylebYCcaKEuFUvMX15tY53MMAPYH2q+o
CTOFcVA60zSwfVEcyRWzVoG4QRxzr4GvdsaAXX1eDw+YoOsIE2ndXM4EKOGHSV53
xaJBWYXbghVCriI51wgmuyBTolkuICu3jLEn2KqjdlanbcqXd0RFYlvcmnum4MFC
asPjrxGM44LUX5YxOLUCg6IkVeGccm80nuMi80LrGuJdG2e5LKNc9kRep8x1LaSy
41p3gzOtA3g501/poYnWm4VbiTB61Lz1nPOobeudE/W9jLUx2W28DaPkbi60uX+U
9wYBQm1X2u2wcneUWXHtQdtHl/tWzYnHGzQiw/1Js7htVbeTO82AUboqHpbT0VQn
V58xmdLpyaekjqzw1zL3drcF1D/WAy+gZ0ZP9x+hw/bnI7lWGWSxs61B412lHURA
qkccEWzlQiPIPniKG/jJW/d1hBMWlPxVn8qcCz8vIJzqCoR+RAxMFGipZQT1zJcy
3vY3vwCDK8C+OuBS+c1X1q/a8IHqlBI5H2K7jF5JSsCf9uf6YokFScZerDd7EkL2
NbTpRsQhBXVkMjJA6qr+k8fASkZW+LB/Tlx8Hf16Z79X5LdA33FMPhoC2oXrckmB
YbYT1KV6idmYpVhg6oQqfB8eqA4f+WY7Mh1iIhnZiTnAmT5Yt7zmkIMynYoUgfrE
fe+6PoqyBK4xvbg66T2TBp+W/ZRRPHCNi3qfrgtXmyuHSGSoaioPB6IBF3qVlOZL
SalFkzMEAkonARxTyQoCbwE7B+WEjprtXt3mFCiqLTCEmyTDn29de5iBhZ7DN5eW
D0/SYI0kYZEnuglNwc/sZGuXNvBZYDRcm4uPkNWoJbfs/1o+CDfDRvQiW+2wF9W2
IRwFS85veT6yGuPEUDBHM6DmEayrRj5lCLH5f5wJxOsC0mfAbya1W9Gs7ijW8jHf
DF6S/H5H5TNW8++0QJPM8MXShivvxvuBA7GSJRP7Dneq/hIq2rFnE/j5fXP3EYqa
NHSMrcH6KsvX7oki6k+CXce5X73ruUnqxyg+lwfnOjryC+bVl+58SnxGglxRAI66
TZs6d3d59vFTXSNCXd3n2EXpKRwGZlZdr+qZ6JL8y8fxaY1V1zVfX7bl5SRBXcWx
HYVn9gkA4L8FeFqeH3CekviHH8ErdtLbtP0UCPqIAvs2E/fgd1mXl9rrbgMY2ghr
tpUIixyxbMo7X8QQMC4rNFTZNvxYxwYEcqDM8pwtAjOQVHdy2+CHNB50txewNYsE
SZ7Byo93PZwoXqyFEOSlOI0O+MwEx8VSH5qSUDDh9xhIW/8haOOXaMExQaZlHxC7
etCZ95rLm9TbcTdI95sezG3Ycj0Qmnh2LzbomlpF78nFYHMwELj/ZqSY0AGidFwW
dExB2rgExdtYOPVytZKd6VCNEYfm7esX0dIlc9URRTVkjTHrr4VVyTGf8v3O6WWv
bYkgz3VdFssiGhTVr3N9liQZndSKpfdxGoy5R+28+9BCcraUveAhzoPjf/inrV29
vbYivOzreWlC/4wl1TmYOAVbpRjoFRXZxXlvJSUAYvjKsZhMlPBPlH4SdY4t95F7
bryisYHhf1LlzVvCZbTo5yHZop8CPfDUIV6NqRLEcj/+H8Q8BgAXLkuw0tlR01CX
lN1ufz7xcl4wwKTjXYbCeMBR4dwvvQpecD2enYORYGgd1Ou0Mp+fy2omCxmRWYGx
ZRuJgZLpiIUITIGgNeDXiA5XFj+qzQDZ1HCgI7oTET35puVWPdiVwV6Te5RwFm9G
e0b2TF4E5fSKQs/5MjIrmD7EijjFFsTD9ZW5g3/jOIqTNVbCbKSWa/Rz8w+cn1eC
YGeFYX2SPdFtunSgZL/MynibN53VlwsHzddJB36tdX7do8+h6FZ0jiL6HFcQXpBF
W54AM61B1JEYqYzdE3gP+4oW1Z7w880Q+fnNnXDvae7hX4otltBPi4mVklfXtS5u
twPtg2RS0ywULSjHnfzsdUudEn7YAe06AqMR24su+JYpb17aFTnsLpW4pdIagtGW
smyfxvE2JcFAIX/x34qy84CNLy7AE6mgLBBlgKfU6SyfkHKwvTnpkStSurvnndtT
/Dj2TatBUNxRI6FMvfEoSzMyL4Btggp5ZM6GiY1j9ucG2DJhlRnmBDMbzNv6/YYV
MEM9OlFqhRGtMQE7uOpiWYG/Dtpq1p7dVyymCyEfr5kQ1k341t6ytATHWl1e+eJ5
dkd0QwsX1RZstL/IpZ30fENd/XDr/4S0vXXsLCaMvcH9438iHRlhG1/8EoP723Si
yDsMcxpqFGWmcNHzNobclSiQ8loK+wR+dHb5fanKx/4fb3EKXfDJmh2UNDIJzLo0
WC18U7HaXUYuuxHsdI7vytkelmXrZ4A8sS/nrwyRNHOV5j+zp5EiW5Yus6vq1j3T
vbvJp9/nv4y1P0hC391aVlSU7OeVCtLFpj5NfJUTuuupKFCvTt1kWjp/7Z6wS3YK
ePTgqm+wE/JI4RDb3IxEZdtxU87HBe/05+GaRmFS8iqlqqLgc2C4xY/4fTzEZ8hc
OhBu/5IbrIRYvWpdY9RFej7KBN8mrAluOaHnk9BWAHmDDYKoWBumyNbqEVcEny+G
rwOUnk+fW7qDb5VEbYM2DtZgIuAfZobJBYLyVwlibZiaoEPxAbbHzESFvWlgcS9g
4bgr5tSsutIdD618gcxKWPBQpuxpablaJUdV9B9xRzIneJVDgc1ufhOweCR9dpFC
SMSWs6EtW4k0p0wOHu0ZfwJooY/rGcZHC0DZISuNQHRoBygFuV0CEwcRx35Fglvr
Bx5et9cm+iXDXsLjhpaQgtnHY56UtEdvFlY0LF5E8WChYne+rd+9QNBpC6yTHPa2
EdTi4JSJ2biy8EIQABExLDUfUxqxw5gccl3tHhcORXgBPS/mrNHudWSgHOjBSInC
+hwAIn75zccpuJStGPe0AZoMn522XCsL6FTA433wnpf8nLmOkSA2coLfkgjKaOjT
izHfjvHvXTE0vPTmkbW1DuukPo41LGDtOAR3NsGTuUhnuDZDdW0Nkwk16rq6MejI
n2vUwY7gN0WH7VErl69fQ7XA/eiu4bPsqmnPobOpJFAEv8ixGQKCWcGcpXRWo4tb
v0UBdrEcXA3aoILnH7bmuzXDu5dXQ8rfJSUMI0Wc6MuZfCy3PnqRAxJaxkr6mVvU
W6SqGZw8d19dt7V1ZhLHJWslki32br0jze++/F9KvTjBqcv9sapiGUgDmqQfh0ij
myq8fqcaOnLpB27Ie4xHR2Yt4wn5QiKevITEGa72AdaGen9PkNhThiSj6WHrG+yS
003/VNOA4lt1+qOCFTCzsK6grkmy+pcZZfAnx4VIwvwAh3Vma8Cv2d0TEqq6oyGK
IEVuK7EszImMQCll7eU3MIZbvQGfK3UDeK4SoMVkDMsQayjfS4EMz8uFdyncHnyB
kLoI8gdrhP6a8BJaRx874w3lETDwK/fc+x8ggPLLCj4nLEQzD2CRGBYGRKp5/N6L
+Ex1+VJGRfb9v30XqgWXPu3ZUjg2w5YL5Vc+bwWyeiXJKSod4OPA0GyMGfCLfsLC
7ExFe9qMp0DBjXXqHt7mJTojv9dVO5h89nNCsM6TQcQSqgm72KZ10XvRXms+WORf
cm4tP/IXjc8zvMAWBfTnvPZ978f+/H+j3vjV/OYXvWqcytvSaKrkvmdVlLm+qHgB
/05mp01x0oEkbH1tJI+DN0JYc2fG6+c9ff+Ctb6XQCa5HxHj1vU3nkR+9cIaT+e+
+qVzOMqxEX8PeK6j9+pam2Bd+QiBYIuF6F1jOn8YKRpO/7dLKsAUtQNDZsR9G9Rl
uAlSdV22mtYW9t6tL7cbDwl3EH2cOJhN9gGv8ravnYnDxA+iqUUqmoVq1ystmBB4
J6ekSSoKAwOFsCx+pSxQ0JAPV+cHkPDIyEL5l9qYj2CDlnLrz0CatTziiy7kXCkn
G9SWSdAOOnu6whg9biEHekiddu0+uilT/Ng379853tVTUg3gFp94YKUZQc/CP08m
BpeXgi2/PmKwatY+vagM7G9ItBXniIkCMg4NUS3LLr0sPLiXVI1JPLt1Zpwftuiv
t8IYZijwGbHcymyWaqU08hbLAQIIUL6p3LreVroEJvqZ9nlIK5y5z7nLUdwTNVlf
7FskjL2UCPxV8lhFb2jHNV0zVrEIUGc4FfXOjOyvVxMZDG/TowVtPwtZoRxCg2GZ
IKyhWKOlYDsaKcb5p5cesd/IimsojNEZShqWtzrm3MFgs0pm2mq5igz0MzZ4Fbjq
iGiKiFjwRhUp8LRRCy/875mh9lqU+h2wDQE9mGnUXJReKQ2KtSRnSxk3IR0zH+DE
wwvmSc9F4YtCWHdc40sv3FEL+L16i3/FfMsT10MEh3urQV0DF2p+JSy6nDuDcDgN
P3BTBJUqbJrEeP9Um6X0lG1ciX7K7ktawTUT5AYqWVUC+5hbN6GD8sCl3vh2pPQ7
W9TC1p3wESaeCjF+VsqBXK4PQnEH7iXc/yMWl4OlKNGJJN+2zGgA7fv4vhOSZopp
FyKf8RrFZNTwxQaNROZ+4a3is8qIS/XsHYi9tC8gxmZHC/tgDxyBBOqJUogBN/y9
IM22VnQfrIWZGxEu56fcl/GzecUP9PBMQE0aWm7oXM412xgw68o79GtL6UTd5NRO
VgXgRuKY7OVpXA3b2TuDzlHdrNzO9AAK5kyLqf309IvpxSXanKAH4JthmOMASz3S
YYZYzITmBPDoKL673JfyCvC9mdKKXMRZ+kjfa52ex0KbuSQrL2eWtFwtkcu/JLgW
SnqdPNfcEtK19PjGgimkETBcDp/VmO4seFsylu5LiyKfOHAGLg0mWBQ92QJSCeVJ
gJfutugGscQga5qCYDNO2COJbypIhLXrS5WgG7pvw7qUrihxeC46DxX/alDe/jzF
18kQ0W1gxQhz6MvfzkGytyvR9SPuBPIc8F/h9DeQFzxZBWzgLyKlS7ykcqVej22i
g3gsr+mBzoy/WiNI/AZBoZsiP/TxFUBYuNrO98v3nzaZbxhoVsg+0+i1fglBlPsE
A29JS/ZgCGDcYTPeqLTFuO/tkXCgw3Uhmg8vRmyl28jJRPRHtjjRx4st6Prhk1Ue
nY5h67KuWvZgi8h8Re7k6xn7mOLZD/KGW6v3NkHh0JiP3ScgVHIlrdnxi9Dd6tPg
r5tAUEcjE9U27Z+1P1cq3bcWIdbnRrFKR0m/hss0PenK1M9HY4XPqjZSVHD3iokn
JAAkzpcMtbRHiA/lmSNOkwLola1cR5Tb7iMdX9kniNfUyCaVxMXaF99Yh6H0ZznC
BQVbQjoAD9d/wOdoRSgBMpwVLJju+D4OBnrtzzNvD7tbYQich84xacyYvV0P3K95
r0sL3L77QJQN3R4tFLUU/eA8lUZGDAI9UiOlbU1xquwJzq8CjgR4EDXNDwMaFfVs
RYoXpm9Yx2I4Gd/ZLdQGVKiXgO1n3VzX4uRFFkOdzTQGN7pxq49jk0hG0GZot9aF
BIMA76peIiMvggJdYcBSloj7w5XClvmS5HlH9kTV5/wkGj4eeA/WZj8byqPrul+d
9acRvEbDst50BNP53yuhcidnrE3sNRhPF3BWTIPvDw8f/xqCjGBnG+9994HPwBUD
9WKVUwHjjccylOSVvx2hjrTvR1j5XI7uonlmzzP3n5ZGqH4I6PmSfSbd5Z6FORyJ
SOUY2WKyFnXFRMBdUAqBfhB+kbvQOzNPOLN8BcZJmbO1+tEF82JVqAMCt76ddb4B
j77vqenB6aNNTiLmOnAABPHzesvHOrDS/f2PrFCt1XryvD/s/rk81OPnqlQAQupD
s98LORmaEFgaxWWd2msPgNXDwRC26ji3vkISRoR0FSgCb/8U36DYXA1/m2B4SkT+
DFcldLBO/RbCZHRRHCRGRK2c6VvhH/3SFWlFHj2jv2/H79GoPAtKPqJu7H7CQ1Ph
niS/iAPvmVJh8Dbb7HQWtnrfvXlIyF6Qyt32qYnXFJEIjzm6QLHgVav1Iq5+5UiQ
iqy/Vh8tGmMi6QVzE0ER2S+LD5CFZc8DkFQCmGqzYbkHoXd8UE8PWHDYq+xc3euy
jTVr8FL01QmjRzV522tzkP2flQIeHGv43OxwqZD/kTtBULMpntZmJZhdovoZ/dIE
1wkKAF5YeL34HTnmZlLbylOe093RSz6sYu4F+YmjmLZebBawCMQFSzlXJFBogl+v
WuXbDgYVIyUON+UFnu0hq6xCsqBZOCLn9OW2wVBZM7l8/nwyoawV2vXJazPTZk8W
PhS1ofZ+LEawDnj/Dl7gAegB2dlzLbZ+vAhX4oGROwarCQtYMPwTfrgvx6xR03IP
J7gWyKUD4Qvir3eVecz2qwo78bf0FLX2VJ/22Lx+abMkqTssacoHOr+YNiD4kvVA
zM7iKf4LU5luTOotiTLBKagU9czHIc1bYmOyGNmzTFe+0pUc4ym/+FEMGd+7kNB5
30IHV+mhGtrZ+kJWzXgzPkqmRnA6TKQfM0pYhDW3524HjwZyGwhyJYIjP8emWG+B
F/RIarPo7sDhdoJtoxSWwshQ13C1tMt2DWPRG3bqnVzOd2/dkD5SW7tYROPH4Z3v
19aKDJ45PJ4mGBsSTk5CtwJyFGUItj/6AeIQdSw/A0+1BDCvG+w/IMlYcjZivOC7
ZIBvqrRVsv+Llgx63YZZ/PZzIVxj5CM9W+3EQHvN4zSnuowxSgZgHijg6Lm7pT9W
vrkgGxj0X41Japv38iJZjPn33PDU/cO/Suxm3pl2n8goW2NSujBgKfPhw9indiX8
A9XjiQmC/6i43P757xNKOvKI41tux+OmbWXzyyild9EiPv48wuLHR5ywhBCAORo/
j0eo19x4+8bGGqXE90nlmYj9EAIU18yICGK8+Ildn0OEXUP4gvEdOZKcjvXklgK4
p1bMDU25XFx8WoQToNFSWFRX4fVVFg7f/SHUQash7SLzVrwGicwl+XKPtU/7wEk7
i30EMmeIEqjUHFCE+9e2eeT88ep+FIKvMy4CUMLFd8QclKTdaL2WHoHKuavPvIqp
4b3bZoP2kcxRPEwTNBNwO+36hf4tNPOj9DUaMQz7RrhokUInr6MrFWS177RXDPlU
dWxb5n0fBOBvDmEWN0c4iC14K9xRN6QDU6MwZuRF936Vglh18OxORdYtubZAm9Qx
4qC0dn0p8b8g0om57HYX5qNgzLrxY4IAHUK3fTJIWPwFk5/k8a0G0/4ySSeLzyWW
TLgc+3041h29TiaAZrm4kJqejTMqs+4MKS0uZbzl9Dly+cOfLb3IBCNPfefmZVVx
5dCa2+iswH9h6euClO+J+576AMUDXJB92Fo5PeXLZ8p+2I/lxwqggqBhJUKA/RjC
PZWfXeteE5LgOZwWEollbaY9n31Y5w9ZEyck5VQu0FW04623Pq1aZ7aFx8qwW0Hq
4B0eXdVlrUacblErOrcNBXWELLcUJRDxqoWOKAeKX8cWeDWAO53t13Xi5z4zNYxv
PfC8V1qbtJctEdk25/oGNm8Iu78yAZEG9ewPQMW2sK8GDNs4OrMwiJq1XwaVDS8k
+mHD/KnblOjTE4WEV7mnsUpoKPE+kcklV2NkP2Yl4eEXklHVVBIpsZ+EVbWVzfwU
brwLMeBRUSvqXFYDh/Dfp3SVv/GSv0AygSRpfpoCK5DNUPsUI+Tu4pO2BZ9qtB/h
Qhm1l6YvHdevvnjf8XscW0EbLomxcQh4s85VJWFeMXG4TBGzlJ5J3exv9CSTXjYU
1p3dA+X5MIDHn8U4mIor4XRVLJz7RFfnGdd/D5tsPLpMAobSHOYFHnRoRTWn9dsU
ohnjecXEkGmQ3xBGPjGNrR33G6B9rPwf5gAs1qGOKfu9NzhsHdpX/OH20TWKHuJJ
g7XgwmVw0YI9YtSu6P14/stRmx0oV9e+5utL3FukGrp+lILSmEuO9osc5+KDiUFl
h4tHzgEn5BqbRjMtcLoU8FMsVHmBFU12sboqkdEez440kKYL7Ex8VNHRCvhFTG+r
qq2JxLLIy8qD8ovKuQFhdPy4TGMD/SK9laQr9/M/i0lVK1MX4YEuyV7Xg/HEH0lh
pmce7PITmEZ++XHY9MITWTeB6vykX0FbxqrrmyI5s5AWKFbn4tZdhhD5jKPWBKha
Og3PnZ9aEeBXPuMcLm/Vtto8rqUJ/kYHzt79z1Ti+0H0HEGvHQQdxioHeBj/yU0s
0IJAsS9kfginuG7o9K+E6ISnlA1+qe7bpAZowID+zwmNdrtZFYJbcLF+j+Oxkbo8
XpvrJF+PMBeKOitz+18n6ddvW7JttWqTDCzjh3d2n4f6RjrxPy7v+O6gC/cbqNCi
DxYKpptCVMRsqL6FP3hAB7Sjgk9Lt7gDrDuE+lBX5wP5zPdL4MCzcxofHJjFkbqa
95lCPwq1JyNw+efutyYcD5VExJph9yI5DjvidomcB8WDko1R1Q2N7rWcD70kov9x
jxD8ibiOlxGEOLjvRyN61it/7ayvtLkzetmtM+qKiygLYjpwnS43c5bsfQh/XwL9
l9QvFBu6rNm04Qxp+Ndebz/a/MjmQpLS/Yvrrb0bN8OL6gKHJQXW7sHPC/PRj2nr
6YmTuEOsx5l/ZZcZ6tlx2DMML7CK48eDOWyml0VYiBb1vjUaXDLAxyY+5ezxjhVM
cyR5/KO0/hobJYHB/xjvGuvKArT0MI3koSeJplF4yLg6Bw4Rag1bHzBVUxClYhng
P8ACYvNm21P9FIEmhdq8dUhvDyVwUc0DO96dgUVbvlnBMSvOQkrK1+upPuqJjcsp
p4Nl0kO6UW/es2KBi707TbHu9eSbDpyHB5o0ctG0YKMe0iTqUTlBTWAnoKxlp/bO
1eHikoYxTUlELS8c2lg/5YE9YMlJYQIJffzRBjgK5dO88ROihSBIG4yFfSCuFbfp
S7dW9BYaUeDaJH3lSiD6zsIAPtBASHlFHxim1WZUtwKJDTMf2B7KwBZ5RiglFIkL
bhwml6JYJyPGPunAtiOG8IYZHWgtbXEN8ENgsC59jHUmBU+pMjWMtKgvZ2+d6kEh
1YFTa22IZdCU0FsfwbNHuWs6FMLEvy/RLwJecFp52dNkjDgzn9NRftYe9VaxrgzJ
RuvqKpfa2qwHw9fY0jhfhEH1UtbVtew8OOF0kALk9dhM2FsM0LjwAb47Ly5IaraM
pAV9oPQ4AnlACapX485WQ5oAlZdSdXaCBrlsgneElv3nr1Cmq65x2JNT04mtYbMR
mJDrjkSO1v0x/er/XI+iPVOdlouvN6JW8yZ/4r696iJT4FqcxPX/0PX7I86M9CNa
ycGS0hXOAKFA7TFqE1f1qz5bMZQatHdzIOnxwm/WqfBSmld7tZbJ6o/iup0uFTkG
LnmMMw0fxnaE/Xwkz4hgXZW1UuyxZSl8wQNbK5FjKzl2DU9md8lRKYg6g+ZjyCqA
zcGpHieiMWzTLLpg3Rm9MQj6TWc4NUoefxCTxv5/616gHh7TKBnbJBFBWmncvXW9
7tZLw1AXmpV87uP0eQ+afFQlhXGALFAB34nkYFyQBnwMYY4GzBmDiI8+qESlHI1n
LwbqQfS4HBzpY/HpoYQnkIAJZiE3Q1I2HtQMN8UU0fcQaooRaVKjr7IUzvLtLINi
abu71HJMnSgRcWkTe40oRubNJfUBuwQ3rZcOAUdYLiCmHw6HzlFf/Izoyvv6xF3w
Ox06iqHeuzOuYgX8Z7M2MJ6xRdbE9SfYTTJ3srAB7r4/SlO9kHoiTTNjvBCXPQ8Z
SaKFVhrfRLbmfG3raheojmb9G0i6tPpTbOWOuCcUAIo/zrw4XBQVc6RINjq5RGX6
Y1QeWYblAkWe95WQb4l6DI4TwI8bhCfF3ScMnUYNkSxVz9gNVhCgwB7Ymk8nu8Ag
rvl9ZVoY9FmvMdxAkH4Wv0g/iQAWNHwS32EnJYjzK+2TjyvwETSKmwOOaUteBQRQ
HkM3wvN2Fuh0Jl3TjCuOF6c/8FSyvguER7GzkEv7PikGy85MfdOWAvazE+kGtdBW
EHjrTbvQV4EMloE42Zj7T6Pz5KIJ8MXGlv9b4cq4/4IetlMK3REnzPzRATjDely6
LY682/Ew5iKjtykm38m11USp3v1zfEdiT0GXf+8TLMOWxFXh821w623HTp4cu+n/
S8fp7jFiTkoJXhgc5HAtF2UXJKQG6cOZ3K9kvsQBC9R2MaSvb29jNiVq8N70NXpd
o8lNA/Kv5Zh2IwNveGnoFPRviPLV69PLCd6MfpHFF9PP0iWceTUO7pJSwIbfv8CZ
zlrtIHYxnU48rBWxMocd2XzHy2QE+Lo8gxmU5vyiuJDHzaaFknlyMdxmu3fDF4iN
CJ+SgzL+Q4E9zKZi3BY6GNYPo8c3JOVrfe9XuFd0b0SrZAkXWynVF+bQl5vIicrW
/VYLPE1pwsN3UUwZceL9KPtxgTkWBhkY2D+V+HGplgzfiOBC/mPVbhZYG63+ziur
BGXEvN1l1ES2f3AX92qre2Hs6K2r2Yh3BntTA7icLDSeX/ReyGuMZDsrQ13LPzcS
akyUfTwwrX+cSggTxApcU7Y6+0bbP6dWHruNPO1F/cmRCxYMDtQDaomvg/5T001D
CadXsp6OKFnOouY0XdOUOBMqJ7kMNtdx74JVNM4nByiqLxYnQ2BNhLja5W9vsVE4
Qej8IhtgsI6Pk4Qc1y5k+ZbVmhqT5sziZb3t5PV7zEdLAM0RO8IjZR8Wk3McyG5k
8Vr8bsI/4u2seSTcaTf74meW8w3U29lvc6SwUL4rHqEa1aSEpV0S6MfrVas18sqe
FiriEXRCbop8ejxshkz8pkMdpqqXiZx9xhRWE2KcimWigxvxLB+1hR0LlFDdZP2m
HUVcOAbUbQ63YNppzI8Y4pIVCwCBWxm+xq2pmHOxXnU1zqJOfx8KHRqLSyyKSKD9
4hzZaGtNQsBTCkFA4TTaoUwlBzlfjDD2/EJiXNF4Z6voYg0EEHjdGc1f3DPdSpIm
0OGfg9np4v8DWoAzvOfSJzdR6Br1RcUNFOwRCvtOdqIplmknwd8oOE7NoN3FEhNQ
gc+YQQipzUmefM+/f8g9qd63lwoKpo8ncZdDsWiDtKu0Fjd4QbHgc9e0AovhCFgz
FcCLOqeY5oHRjybAQ+UiQrYw+BVlBp9QC+0ZhrvCD8DOoVUlEr1lKpnnHJpatUOz
XMTAc2stUSKUKF8eHEHMDJkrOqFGD1nX/LFowaudg2++1XSN/7QBzZJT6oP5aKgm
ZCB6OhQ3bG43KqTxIxmj37GSDKPuEzswqVXxFsAjxYuLawjrDp6eSv47gsOYAevT
uwh26mtb15+O7Ze8/P0LGjlmNDtjnOig+rog+8WcV3BAVH5Y+/a3rYXE7QlLTbWe
o2VyricOm7YYU+zM+x5aYwM4neZ/Q8/L94prxiy7IkzQJzqlx9E+YK/K4p2V3OtR
oBV/Txbr4WDfnveX7pvKyLLAsRDRFj9bp8ZCESnXkMcKXGbd04hlK+5RTO+YO6kl
Ab4C8abUkuSixSHZFMFbD2Ts/+CM4FFNoYmtLaK4bvkWxfr+q1qMe0MAojhdncIm
Htl+5enXVulgujPceExHvWH+Uu7fqUuSdaCwImRcj5TlaB5FByEkSJlQWJYpe/A6
Ei3IvxRLhhmSvaTPHxRCw1q3+HCouseWyiLrLJ1Zp4zr/V5SqJQqSNISN/LawQEs
Q66hRxYnF0GJRXgGtMNPFVrlA5R0uwFJwLRKIGSlb6tsuHpG1onDGPCOK/sR3FmW
AXNXsd5uz+9BlaQcklx2+vFLEYSt1YeCy8oHHAU2fVWCLO648xp1TDtArwBGxfrB
qOC0FufE5oomD2HOp/MKPewpxnFPB9u5ITQswuk1RDvSQ+GRLxITdJBw35po/y20
qBz9QyDG7cK6PzjfKQRV066DGvZ0u6rykgr19hfzCfVuRrHB1S1ncadoQrZNcFbM
Vpa5v4dLeaBWsQUxDLj2YQO3g3Nz0qhJrAzOhbzC5hC7MIFEw5PUXd6GoVsH0Kv3
N4vhzNHzi0R/VIBuwhaVak152PGWV8jezonwuRhQT1OmOyTg5rHAJex/jl1sVPRN
C87xw7IX3GMlPsYyTQjYumCAd6zZuewgoV9KngacHZ/hyPnFX9iaUgiZhU+fo3X4
HaVi19EHdRtTmWfxXLMx3lAI4wonYLd7y6hJEm/zCmoaPdFonS5VEyDgHhg1C5Cq
2g05LAxQaratyCnnCqKioUU9Ma0OxQIQaClTMmDMwlHa5xux6pOqrkvmMc4Fa8ui
M/y71yMo3kncIflSp0ZBXFfiREYIsE+FLC1AcBpsuHTxI4uKTlcvrV2bc0Lpu0ED
hXM50sWsMzUWeGemTh4e0MsP/I6e6HiVepeZFscRewL0/gOZ2hMVndhC4GmjbmFA
S2LDkaMmZ1AdEN94V9rrTTxfbWljMfpY1th45gK8ezh5y4LqDwRnRuxW2WMXKwqy
TbWcVjqf5AKuGqen1h2xrRBx16WNlu+cyphYYLftCJlGsbKy2iHSgoL0I5/2iJBQ
Mq4fkgPbQZNgy93RMbxiVL0J5R+2rO3JKFSTubBkGzgany1zMkfMtFSOM7npAWc/
zskV3scBSw8gmmuaIZv/r0e2tDHJ4cqlNzKWKBlnMiya//qqyzLRt2Pl5xrs8P8b
xshyWM3vYwoyI7WqCrpvSxGuszyT5csVHm45Wq3jDCmgzgMIVLyexBD8w+HrI8MP
8vqE1n/TwsPg9h+Tmx2Nnn9NnboGDX6ZT1lBFbe1jUUwj6IAxrnJGS9adRRF2uq8
lqAV0T5WE+H1+LQTNwcoU/lV3WH+DFWAPj4UFHW1rWi2HEnikgHOs2ilRHYwSWEd
iE5DFHwHBSghD2rL9BavdqWw0jX2hIbHpoYzG83NeNaOqRdYiU2Mfn1o2JKhP06c
f9SP9VxqJ1daK2vciN+6bw3eRDZjdbIoZk+L74O5qvJumujCbU13rP5Ss3Xs6e5Y
5MUP8krK5NbmzJTT9kLTk3uPa5HOlxme3wi9psbLYMhOXSvxsf/73b/rVFWFK4fV
xSUR6kFb7XE/fg7I/OzCYFbV1SC9qjsvAiMCTEN64aUaq3O0UnkznUDpCA4eIGTh
CqkHXZeoegqhaHmYgw3j46uvPx8Bu/K9ZJEaRIhu2VsHe/l5bUIvrJRAZA89mrlc
7XI6XgDYFWlTD1WbsZzo3a4dItHSjIR2aZEEE7z7mjBxbKKsJFWzKruCJkvqM2ix
JUJhDt9/OUPPvbuQ2XBxUq2kDlMltzYeuomTzpBtIPNNyQdxaoZe/1wO7r38gJGj
CGyjsleSpwa8jOKTlsi8LtNOjHrTCrk4ycqNCQ4j1OpNwri5PepwdfQC5Zc9O7LQ
z3GVaUyLTTC4CPxpKIOp8ShewEErUdPHVSkUkh2dtC8sZPZHbiSW3Kkszk+3cnjQ
Zr2IRzQ7wBXazWhe16XHuv+n6StwDqc6m02XwBalePxmYYWXTmUo2e/jIEg3jaN0
B9cWzlyJT36syJZhGjvuR+u+EynGHPov69nA1nOhMRIphXvvXSgZzM1oNJMDQ0Yj
XlAwPusUOL09CnnD1VxxELVCAk6g1bETRcnvWoPvciY/YjFMzLd6sSztlJseT+nV
r+q/bcUxio3pOoJfqZ+AKppAXPC4Rzh5M9WoE7fpsORT4MpS1TbDn9tZ7lRi5I5c
+fgmQUWcPvRq6evEqLQoK0JF5XfVJuM8mRIAbQiFMgl/91AZIdSTM3DgQtqWdRvk
MC0gIFXCRMdFkCeYZLucZYEeBd7Zf3bHzGOLxcj9IKDOyi1XxnKTu0g/Q+6FWMfW
Jpu8qDa1P1W85pw8Kwccd0Q0jZwKypPrmYPmZt9+7IQpG8bfhi9CfsZOMtNnwI+n
ZtpxFh2Pt8cMa35lDR5XRgHTSBPeobK4EgsMj3WxB372bB6IW8CneRPt4y6mrqIT
+GcQgpWK4Rf6QsLZ9IZjNMXkDgVOMmMiaxLgxgaF7C8UZM7oBBls9WJcs4yV9AgM
lWr0V8SGZZ465k+zVpJ+E1fnRQRdeQsF7G6nF+xOt4V7EUGanaLn+ucK8nHyzM0P
bVg/Udp5GVz/nBbgJwlhEWD4oAc/ZeQmzWRPcIF7YfaVv7vJRbNIahzUrkD35oZC
uoJksv/n9ZMM34UQf2u91dwH35T4kW4QWvz7Ho4bbnmpphDnxOSrsge975cnGBiz
wgkfy27hnV7sbKYoX7z+bTqv8H8Ex1q3Jb5g/IPQgkdpv4KF9Oe41P0xPCyBNt7V
hEVAuG/22cZgHAR+VS0thLku+GUGBNfdqbk3qRFZbSCIuCywjlmhKKpKcyo+8ibf
Ha/OE066NqTieKi8wZsTzcddaejoXLomtPlxk5jypHCtbWnjq003aJGUX64tniIG
PwYpPOzgihh1gcEt1hQrYFf90T61tRoAd8g5tNH5TfByqT6REzPc+zNtfS4E21qI
uwW1n26pzEo0ZUcoFC+movB/h+6GJYiyXxAUg9ySZKRmAuBaY/T2WRPj3x0hyWZp
yuo8/ZgazMUvNUlkUvBe6jZSsa/om0HFnuNpYUM4HRIySvDrscQ/pHbI15lZMxTj
5SRfUchr1wASVi9+kLsVUvJbcpCWSaGKruC5weO3O5winv0vxkkpYXHd1xQtts9r
PYaURbj+Pm4jc0PNUbo9uKN1pelFNaukbev5F3n3yZQP94IFwNrbNdYuhtRk3jY2
mr8amXehG9F1v9D3XooOGKKrJfulpQRaBbv6eLoIkP9JR5UvwEPFDUnzHvTOGByz
yn27DhLYMB/Lo7OLtv4DkZ2j0Tz72/TAy33abrdEHzk4Ym5zdm9/kPtm+YWrwlXm
fvqfK7vabdo8nf5j+2hL3MNc/2AuLv7aeZ7zM94Tfo+8PDVWR1iudIChc1OJ9w07
36RArjm+2hn7mCngF8dWTGD+q1hnJT8+f+FX1tL90mGZh/VjXzVciijrAbPFpJOz
RfgCM4pHvStLJEhIKO9Fy2z9yZzrNammA+8vpOrSUE59TyFY7F6q8cOf1Ybbrxux
EpXSa8mhTeUoCOlxWVDrjnIQIiJqCEyoCn2iNTlsglcLHV4MpJH2Ultsi6au0n3e
ihgBwHKpjkpFbmZxssZBj6aeDp4lD02DewzQH3wU2TEB/0oRsnvjJ6pcNbIZ3tTR
qARctY+FegyVtCROjuPRKc7lgXuO41xQsa4dXFgcx9EN2lC8wLJDN9GIWHcUiYO3
CFkNJoETh2djRZ/50PhmczTknfmjBr9o4x0m2lckik1ml52bHJnJmZ9gdbMk8PMZ
dGd8GkCe5dM/2DvLEsVE612sn3eaBr0cie4tNoMSzbeRj9baZm45BMqoLzFIQUc4
oKl6JuQ425GDbkRVSjw6DcasrfT/7CFFfVRISX5ey1c8wSHCbfJy+sefOEMO5Mkt
JOEg1As+gFwZWi1Fx2I/zM0HjpB/c0UhZrQ7SFYyNRZalX2UgCqL7/WgKWEq580s
XsnqoXgMGHZI1Ok5Hd6I/0vqJCRVe4jK2FPO/fVYW3B/5W/z0gf6WCJeW7K6hSNY
ScoCUolgHA7/Enz+URotTqHybFbAsKBWZmBnhcQ2Y4kbTOzea4DAzL+YCUW8x3HD
ATq1h5v92XQMRgsBzBJzxQasKg10z+N3KlYsnH2olf5q7CXsh+oP31KPc+rsNH3M
q+jz35kZv7QLRLvAHFgIM4vrGWYTg73efjpRM8EIk4/OV4ubfq06rvyO+Kxv8zMr
+a/7d5M6kQM/mmqX/JbDznkW5OBJwSOWy+9zpHX0mWS968ij4Spgd8YIOo1/Bc3o
92EnO7ulTPTHUYZEMOI5qNf/mjMYeStDTHwUnVFZLD/zYlPkXt1IwApHWrUbCxmH
/QQA6FwLPlQk0t/ie3fauU95MAwPwrt+GCnLjXAgonODBJLmrwnDjq7sPVQIrEX8
7IkPRCO5Z0tyD6UNI4eBsrOYXm6bMX2TwP/vIfVI5VsMcXerG8Oj6IfpuH89K7LF
E1GEiYkQ7PFHM7G4H10qO6UoFSEL2IH7LTv+C0VaI8z5TgywrxII/8znOYumY9gi
JnDhFBK+5dXSNBYWzLwn9INWhSFv+2o6ntEJWNyAn41ektZZ8ZUlkJh5uml4Y4e3
2jyd/OdRLpzCgvp9tESNDhcigsY2ASm9jVB+ntGNjJl54SVm7pnnyg66QdpA4Qsb
JuYITvE0t9dxbjI2ZJH83EkJ0/OtKBhmIKxi8IeEv6GIekQ0H7cxwZTr6Y/Wupuu
yVFMCV5UTKKGe2fjXTaeklIi/acdBs17caKDmLMO+9Wwz1m50xoBOR0PukisV1Yr
rPHOYerDFIq8db98Jm++tCKvF3c1a/QB5MVqZqGuHVr4Guwj5NyayJtCuPhZia2D
/qj0prbZDowMYCO+Mh/7zG72nOmL/EqY9xIdSPmwnSYlGmxd7riqt6uoB9aSgNPT
8Tf/7P4pjm7Y0BZ7iCraICg2diAYcArdQ9mzOEOvcss7u1RGbPIJuWgVZE2DubKi
76VE/J9A8394YsdN0DXOAZF4sZwSIeWXhW940g681wiTsgK5iRFbG+1tNB/wFFUm
8zzVgpN0ad0r/1nDaNyXB2YnQ99jL8JZ9PSoDZKkSOz84oZwyBg0ABB/auElLyWx
9nBiCdS+88H518QldIeQgd/7DemyN2iLwrNJW40I1FLkva0SkHZ5DFVkjhVKoCVZ
59+AZCAyOpO/DeeqKnFHtqkvS7pPxfNU9Dcx+3ea0DXkCyXA8Bmdr1zNsSSNJ5m3
CdWNSXaxj4XLNXQaEVUgk+gUkFUrg4Xh7KKd6lusyldrJDsCOrtLLs/8zajCYF2X
jxLlbfWdd1LVexDa2ZegRQHNOoGrOWV4nI+Mcb0rs2MUNK2SKJwWRdw3VDUPIz98
cX+M8PqSdwGlu6c/AUoqluL9FNZPZ3synEHD5mm6XDAM9NHLSLnHjipIvoNO3p5G
UuadDr8DUfGl7QUUno+LL8Yepqd89S56onOM70vkid7zet60ke8gPNzNROD3gWqG
cLZfyD1S4roLitfSGbkcr4TLPJFcpqOyknsIYPsuZZBgacV5yMul6lRZRlHG4byF
52MsEauY1wBIJWMAkcuMwYsiRAIfRxJ15uadw7upBbuSNXN4RbqzxK4eDkWgzSSj
x7CeF5MzrG/wjPki2tMohRnwLl1w9U5nDw2jCHQCIh0id0UXc1SRWCbtAgGeUfPV
ta5OdiWtyMUv1lcUgQkW0PUBmMRs1Xuv13uH6Ku42764UIVplMuBqplthhPb2Y4M
ZOxJpS6ueDp0gDE+q/+2APNyp9L0yvg2v/U2S8N/WP4T3mHOoNC3GApHkmh2Vggc
XNhwqOsHPwL+tezxqyY7r1MxzLnWSzcBFKW/5eOazwVSWNRaG2AAd7xouV/T5c2L
xn6N7EIBgRw9Za60EiMSPfpwoRuPb7FxY/zBo6jE7DKNiXFu4pgi61r+584kFIy0
OhHdQlb5VClNpbGBI7TI1hGWVKb5fHdrOOmcx+4xyTGPcEc/CwA+VF5PVr988B/T
xSlFMtwvIxcoa2WVw7kpNaYqCWQJ/UMmtdH6QA84j70QQ+z3CDDvTd1AGv7x8Ivq
j+wf492BpRxeUc38FFYtBUAGTvCRuLI57MeBBCsvL33yluY2qokl6iLsGI3KgH7D
jIfOibDn+jVIDfwPvFHvILo46EKTyMPjz/SOVASurUI1uqHdqRnb+m/d4oJuqtVy
nNgm7gGo4gKqUc/8+m2jqjh2mnr+z386KoOzWL5BvRNvhE0S5xECahfTz6G+0rzp
TrHBNArCg9lztzPgq/jLEWdkjrjzv3v0N2i93IRL+qicEVkGKVo5/6dXBC3gBM/U
4R76A0w+rZrv24CXfusbtVEvU17kzkG5By/x/qrLXUd5I/djYNxe1895Q0IlIb+k
W0qrBAVaS2mWQ4UwfoD792LAyXJp6QCFnZRaBcOZqP4aFZy6Cj543BH5IxWnEFvQ
K3L8/LZzCgaOr2Fa2R+9QEwk1zKVa1oAfMkSSv6X9sHjmnU8HBfiSnYOHXWGtAjh
aYCp8Iv/hlzB1GD4l5ZLS33Dxr9GGAK26Ln2r3EPNhMOUkU+dzNbp5V5Im1XfhhV
VTcfJh2FBgalUxC46l2MTFhHShPewxX2JXN2tMUWGwFKwNf9QHTKxdJ8IsobWuvd
J4/vu/oEbHCj8qcgQzF1OGFW9Os58m5spde/1vnQg0WESnwL3A4Wr143HkyfSEn/
DDZAYy5D//5MzAqszBi4Z5hEUU2yObKi9JfC1Ei4Iusg6gp14KhaB7ocEZcBlUwX
QGOyI7xhHqyhepi0GYBMt474RqF5x0MsbzOoVraxw+i1bbGZNcxGGxUNGDE+NF3Y
9Cu2hW46M+cXmERtl4OqBU2OKPUOKnwSJ3iWyQvbJ8TTPgFKiBUfX37e8wPdeosU
4mDbgYky55J15YzPCOC1Rvh1GdsBlwd5hq92WaGziRS+j9QruFxy6q+ZIIOBrNU7
N9unAHAU3NMqFUj+8ioe3/sO+etX1WYVSF0JH4sSQgwL/snqd+t8ZhrONFIXvRGm
2t1VWYdEyHbcfv3U29tjmM4ffP/TPI5KAHIoUlEI7QKENYjpCuSPi1ngu71WyTgZ
iEYQTpdV7989LEsAqc5wlK6BSUyyQ6fX300LCPiKxU160M5+I5raWUx7zk5iASa8
e9WdPe3hjBDWCgxT5QUy65N4UytFaOxm/cmrqvdbuHlAS4PSd4bEUu1G/AzlHWwe
Q/M8GcubikYwD2RNCAUsy5/zgHZc/MyywO8TXGAVfydgtPRG7qYl/ItQQM59yxuB
WQj+nePMARSgZXlpsJI74rL8fRZ6d4uf621ok1AFEPrMoZ6ATAiRo+3AY8LE+ua4
9Y9iQDlsyMgJ2j2EVnLrghvDVfbbSgXsGE09DIyym19tYW2YPPvVEx8Oz2r/lBEx
C9uMkLNEe7mdCvI8lSal8TxSOvpj1Lffsuj/JSPvBRLhIs+aRiUlUSdOoRuY0up3
l8KjOV8QBklSDx7XaHw+ZOCqY5wqTGSPxxN8YM97ZntT+38aYy5/z5IB9WEj/tWi
VWv94lCrTdRjjvqtDpe222pgKAWBmqklo6KkdbqOSrXO7IAiG1o3AVM7d3vsCNYb
99aghHOGmHXh3C2NeSE52m4a1CnCG5fUwbu2dxaeAChEqCnBZKQsqJ+k6O+tQEUa
pSC+bSF4WisRoPZyHmIefJUkFxZnhCUfw0j9xDCl1RI/yUdj5bj64atYbYzzFjw5
z/1sic1ljgQS9hUhPMbWEMsstxY3CY4PrfKFIn0iFFTcKfyON/HgR4mfJZv5khVn
XGsFrCg3Kc/VuI/wyiGU+REqIilMqW5C/K6hB+xJ8dy5U9RbF1QyozQdee3BSlKg
gOlesX6mCcfpmp4PhWqIdcSdGt7QJMV6RyOPQ4+koNVIHEmJ3Fwc0mAziCfoxk4v
2zpzRom2c+GPTDzmf0rqHrU/+IIfMRND/oiWasQjg3XGqPSnx11uVzXwJDYeh5Dn
nf9vTDZPcNO7VChnTy6XbAJkzL54JNOt2S4KM9oIYjXIDrtvv0+aruQJgag4dNww
jIoI8ZaMD1tdk3h1bK/jTqqpONMQJ46eoVM5857ysF4=
//pragma protect end_data_block
//pragma protect digest_block
4cesQtYV/7vvpg4CBbH2NTV+v8o=
//pragma protect end_digest_block
//pragma protect end_protected
