//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FmOWmhDJF/pMh2Bf3L/vpRsaYY4scE0f+bn+shuKwQkPVhYr98XLwSG0anEBQ5da
T4h7dDn8Mio5eBfNKTSJxSQoYmmXlBS4fBA7XKCENZfwrkyHZ6UMzu9QUXr0tth/
KpGNHtk9tVzE9mU9k3/nvXKc8516B5SEyUEFMSxcGxmQp13tup4F2g==
//pragma protect end_key_block
//pragma protect digest_block
L87BtjddpAfYr5DBp85po4IbFoY=
//pragma protect end_digest_block
//pragma protect data_block
FH3ymjxXdNbWlztJwt0IzBRFOSu+S/AWgULRpi7nayW/MI9dg3fpwikoWnTYfzIq
qviGeqoFNjza24VL583crM3/39Vtr4Il2g1EemJS1eMXlHvRup5KwxuCwMeDZbR8
Rz24UqyqwFDi9YAv7Obh1KPuk5sCKLqe781VMz6MDtlmBoJtkX80HphNYLBBi35q
mzX3CnNV2feiLa4tgVff9d8NeB4jrWDZeUEDGBt2BO5T4b5m8lOgSCWgr5tPbmSo
rBCn+bWwvYvnbCm728l60Kz3ev2aWR/P33qp/7Feco4u4capWzV1y+OZmNFUHnoR
j5Xzao9xd9cZVAS+f/8eYg==
//pragma protect end_data_block
//pragma protect digest_block
JHuPwnnrBgWYkJ4MC9XqyW/ySHw=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Mqc2WxQA5xsaWMxG/xNmpeUJWEll8O+0jCN5r2/hbPE3f+1SVSKr+14u89WKKXvG
dLZhiMMdoYle1dWVlCIMnM3YkB87T/2ZgCUGSTkie9eOJDj8GEdGVcFB6jKIat/r
nvYXyic6+9zRqGWxuneb/TkOwue+7yhRLA5FfTAhW3YMr91xvTgLcA==
//pragma protect end_key_block
//pragma protect digest_block
NWWL7RZjBbjd5HWlQijuvawIdfI=
//pragma protect end_digest_block
//pragma protect data_block
ytgtl4cY8dP0LbYZMEwx+HFXLPDDOiC5TNU6T7gLJKVD426kb1gnCyQAz+WL3CYl
rQ8NgGwEg/90AYejVJF/BfeqSMkxuCbo95ZYWyqx3/rn/opM3/2wSwAILKaR90KO
G3TmrqTnZiE0UAmMz5tYr+5UyJL1bB9UvuA5BDNWigYE5RzjXJyLgIXEYrWKJeRl
7zpOyMe7VjYeq/BDnJQYFumVF9uRWqz1Uk01k75TlroBXxzOfST0WTY/Ylelk2fK
b0Moefb70D0SzStDJwomECMOTmdmtLPHoMy2od+ArwzW1VnCWQbKiTZiQeWx8NN1
2mO4Z7zjp582/3V1hrX/tw==
//pragma protect end_data_block
//pragma protect digest_block
pJWep1Qr7ddYFrNSb2pqtYQnfZQ=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/tI5hZ41CtsmCGFI4pZMhABJEemOcLRStnpX0exH+F2IPnnwQ97pSAMMkEBG4oLK
JC9ND774t5lr/x0WGuZY5pjpBDd+gcQ2qqQKs256Ym4Asrk0LaYic+TeMNg7YN67
NVw7pWzVIy036NpSHoJcbDLhhK4xzYUNWyJkjw68dH6sArhQ14yw8g==
//pragma protect end_key_block
//pragma protect digest_block
D5xnDsS3jSETJabtVwmF1ErzvTA=
//pragma protect end_digest_block
//pragma protect data_block
kbrBw7pvoxxZPvKZ/twyiOVLEtyP8JTNpGDVqYFO3aR5MQK2Mu5CnGu6ZtCIyeO+
EW0tZVX7dofq0L5EgiGQVRgolpfK+oY/rBqsZw//Yl68XjLdvNb3xLeNg7ItTK03
+GSbS7CNUIc/9lY61t/YfBjyuLcfcJKO77D8yEfyF3PTkb1L9o1qHHYYaedKL2bW
TBV54qDFEk5yxviuzlv5ZTerEHFMJP2/sDSQ94hRrIxTiUiCSTW/yp/xHhmtASUq
epLgFKce1nkXAC+EJrjBpbrKuZ20gsqc0dMUAnqm0ipWXWNJphtcXLDwpNDkcZPC
S25zf0exmVk2QkWfBmqhnEDGGzgOQndVOj3r/2MQE9LPk+9LNoCnMeuffXoq7fR7
204EVJC+kVOyUq5JW1sYgSSl/NYqxhbzyauKG3YJDP6i8LG2gg77Mpk6hJA9bZsg
13ISBqDS2yd1Dyecax1vMsA3lFnwtly47E0xU503RvivfYtmju+Vv0Chk2UO+aKz
rZn5vwZCBK1YE8/dDBVg9dRjzfsgh1M9pfNR2hxNI4/XbEUTa2l1PRpDiFHLMY19
wR2W6jpQIVHSl4U/nJJjy8g9425RFEj4neks7GEKWd619nrRQKAVogTIbvdwurUs
7bu23HuylVjXCYAu5LgAUK3EOVTSMTyXPK661Vt+uc7tLrPBVhWyoyqqmm+pi2ry
E7V2KcchTOXHNZSclu58GdkT6wdW8+cMnswQXaE8vGWhGZyAaj2zPhx8Km2XCKzT
K7vRPfLnMZKc5JT6O6lUmp/u/b5FtIiWrTjEPnWSUohwxIymtRMbO1T7g84eJvIU
54GkVGg1PU7x/98+T+qsOIDDWxr6ZBLjKAMZEKFz6jlVrVTBOV6M9/zhuwZv2r/u
R37mC5IBjQQ0GiTsD6Wp+4uLla0P6fK1CThBG/aL6nwIjq1JEusd5apyQjhRHmi0
C9p8d2MwMil/95ax1bUc+wUIZelbmuLYYxBf9hvDeEXEOV+nxxxyf/L6G9PxNBU2
TeSobkzBXKk46B/+ficnbDaTk93pQs/G/wAH5VFW2zIpJq5p9LErg7uHv6sxxWNa
qrVBDzy0emD52+RJma6IW1mrnL0NCTgCUvVTBZoTQU1lRIRfYVnP26jIH5Us9Z+h
v6rSUbzd2RsnzF1XVT7aEIErNBCik6K9X5pAQ13722UX5WXBq7BN/4celepv90DJ
l7/Z3RPt1jdK++kq+xIGX1s+ViGQkXFs2PWcQXwa5jr5dDLbezQbmktKKSh0Ur2z
qW58AvqWdqqUnafDhfm7er9nnMS9FJ71U5NjG7Jj0Q1eYCyWq3WJodV6QPim7rrw
BV9FYmSR2soI4TgXGwfn2QgN0v0vVtApkqIWqfhEJcxLOWvHSmNKmnIms4njhygz
fAUgFqqlPFq38IWeJwdsf/ZoE3Nppd8ipprV2UbO4uop2Uxo1QtRIRivHigyZF8W
M5LPef+E34qLdJ6+sj7SOw7nKQK/SxGjrA4yhG2IPQATlptte52QJb08dxjmhRQn
jRqhK7BBO1dtcQHb7Eys+nNc5ZLPlOhrZAWFWubCn29chOrnrii9Cu85G0TLcSwR
0ttQO4AnAJcYdUKPaV7RZmxJ08C5hirQwAtKCRd6LD+l6hQe1GevMcfk7M00hJKa
fMOB1TEpu8hfPwQBg4ZtIQy16XrmR33LkvI6p37MZupzL1f2iF53e3EhNq1T2zBW
QSZFfgUfqGT5kMekbM9619csfU/uVgfEGiDqqwKTBbH4uITw8uh7BwT7+AvBZ8qM
rzRHyFDqA/NT6JJYw21avESmBd477eINEGpImls60EPo7H7Xl9IwZy8a5aYnwOiE
J+Vi472T5gWdGGse3bngxCY8FyqjfuK3qHI36WLIWDSPd6O0HUkqGOIH0moaWamb
t67Scgazr8+gtL82kQ8HuvCVb/o7SWlT1+Eyq3YU34KFZm3924HEqOuuO8NuKMSG
I8qch+Yzqcxt2sAnEsDBCP0QG1Wwld9lOnNYd75E+o+8W1in2GB9a2mosWirH5HI
pwIoV5Ikbfo2e1PV5DuQlstiy3ckkz+porOIUoPTb5aHaBSKJpmLd6ymFKufkyXt
Aygjc1ykjOT155XAeqYzD1mnn6Mk/e8TuS52BieJNk5tUVCKM06PMR+jv5BXP6Yi
PEr4aGPWWYCaPHHa7FKzMcLcGSHfdFazvqVtCnDdHNlAdK7Rd5xhsqYn46qNzk2O
AqRAMaLHSabMedeMvBHKRT6oDrrJjjKOsTpYuW7HqM55rLqfPHtOWvUOm1Z4lKIn
Z9a7Xn7TZlqfkiHPpiJGf1bmOuI46q6Z63Uik9wuysnQ4okD+7424TgwqGj+vYD9
n87CMllMUmxk4+i0tJ2x0WxAH1o87xYK8gaNjwcKwivLQnIGVkWtQhhU7dWGOcTI
cV2q925jxVFLGMz8B+RRFra5aGg9TbdhDjMZe2GBfSDOhvfgpot05c1ja2XxMyDb
yOI8kT2rAATFt2tDKB8avP+AhlGLNm0EFHZfknwxbLBy7zODgAcj2bqKObOzyyGW
yXZUQMVCUK6RqllfSA6vO92iR81pioFUEqynhKuRSaXNV5TX4dTBqgExR7Ayun5C
vnJobAqmm7c1kM8IRy8/Q8mgl+ZF7NT5UrJy3+kNsimff0/Ca2TjhEWJV1IrfXq8
7GhhiULmD/Uz5yDuiwIxcYci8LUw/lU+5WjCzPyQzyVNLicBjrPD9lI2g5LQX8QA
zuMaFjLnaNSY1U/793dn9p/K6G86liMb2p9pdo+R0dgSv9wdeSakAMIxmnWN7vJJ
iOGqk2uvVC/KYxpsvIMf/dpckTrjuwzpGJGGg38M+mWfHA+mL6uHn/tGOSJ0tWmH
BWwXRFNTrMPB0PR2yQlZop7EeOpB2ISALJEwuBUDSFMTDkuAimHjPZ7cGAiGhJiN
6barQZ9A92+A0ZFVIKO1iL/vSVfK5nc+EOney98NpoxX2NB+W31YJ6RGae1BEzkg
SqKHIotx/Ls5XKpNsMCuArKaAFiaokKcins6a4FJfurS6Y/x1UyhihPpj3V5CBsK
bO3Rn81NjqiRPPOyG5vSLfx+78FnlZyoXpa9Fo7GE7wbsZREnX1SujQE0xl76I2X
WjP+jjGc4bP8bcpr2A7jYk5Q/q1ZD1aek1VQDk2+RwObPhGHbm5Niy30S6hVIy8h
h/6qZSP4MVsQpLL1tS1ybSHVv0sPrRT+QUF/5JrzsOS3HPTd1stac7lCzdfLzeIU
1sebfq0J0xybHSBLHN955Li4dk8Nwnx1U4g75dWlIyOyjnG9qJcpkuc5GLn8ySqL
ubt5zOQ8NTy4LZkrDtL3b1uuyEjzgutZ4j4dHPjzA9GQbR2SgkRqfE2UTYFyZgRf
S81ZquwFkqTSODJjVvW+ROSNZqzLpVWv+aFi83DUB5lersViEhrMYCmofncU+uEQ
uCc8je4ZFJ98vVJZHqbtf8Wk9wZHSkXmuDZsl72h9YPMNaDGyfBGipzfG0C7i1yQ
3M8lwx34kVory3Osv06sYkxDCFLigyNKodxF3A02ugNk1zXn0VV96xF7jrIlJEdl
v+9H5KZ6bK7Fx047cqUZLT1UgS9siT4sBCMxKvfKDSD1nsF/71JrFWSBchbaJxDg
745m8OMcdUiCISqHhuW5wtTij2u6z/xqgW54IdWSsSSMzgtLtOAfH7VBFjEZGZKS
X4P3iBxWkdm1g1+FVGpl8sTVAn26zMekYpUmCJrVT6H7xUCMZT+/QXrc2TMoqoF9
zOR5vosaGqRbSlgMm/TICb4BOazKyAF60y3IcgP52OPEXpWJCZpfVhKuNE0OL2Fv
6FFpLJ2El9a2xMJuf/vmEuFK01OOz5vjlqVjU8IGcc12f3r47bb5jZwjXmXmB3Iw
2mJYY62SMwapSn4Aa6ylutE5R0+QRJO3AiymqD3B6NiO49qSYk3xjWDGXzNj9na3
YAqKbIkANYrfCETixZOFRG2JJWHtCvPG7ktKv3mcyCT+NgWCATSZRIlVXMm9XNk+
0JDWaPESDyjrLcO5OFtIVjAJfTQjLnbYkDcl5MzY8Mdh/6fX42ZAfn1BpoXG1qgf
SmpOGxkLAJpFJSYA+cxgBur2HRBHzLZlEVrsfeViPqWi1Rg30lZ1AMtICQAVk3uT
EVAxPy5L/eNeP91J9ps+35nB7UYzSxmta5/etc6vLBlOQ2f9cyW/9j2fRu1gUytr
WK1cuI4+nut3GpmKUC/4SWJsju06gOQGgfpWpjao3yBcUfV9qlmn3i8OiqZy8UR2
/DuwDB3nNdIcfehegjbC37SXvyMnHbncFXAz9WzqKyuNpjwNgafoSGNlxrfhZxQf
HljZ3lZnN3/uBivfdQW+yFn+UjkadLDkwM++DZW3qE0JYhnHXLn481AUZ1+vweAk
fgrg1K4CdTA1HVbs18aaD7Bo7wRZYmlEOOqZJaPLPghs5+smtPwrEdbCNApm9lAO
S8QMKLslsWumyCDoGT3R4gcVPiKaSi5CjmzUgSSHo5KoQZE/Gjgp1gPkliufP8fF
ccU+VrNjtPFwrP41c+hknueMnNRqeFxKiO+oYlEa0DmxexHjDAAINvqkAXLw20cy
6yorrcJeZYAKLeSwbdEIOtW0iZrS9DlCD/DcvQpVPuhoddvL5yP+B9sv3EFo5B7V
+omBGScjTne970IfYeRnsIaOOwWEAy+ahgzv3j2PYeyICUKFR80FYM1TKutwR8Fp
oy3tM2FmZTORAl7MMNkWuDnfmNuT1EC6acwGYG3kr6WVjx6JWkBk2Ykwa+kKu/G1
ji/Ontb/CHAOM0A20ttwmNw3AjJ047R3oayVpkKX0H5COPHcOM8jhwJ6GpmtGTFs
2HJ2gKPLU1kK/DevFG4GUmjG+a8Zo6VJL/Q4znKNXupDiZtbquWj7f6P8SzrMIym
+UdZaYylffkw3otutoMMObnGIU+2th35wRFmcFJA4g7ICns6DRrieFzEWdXiQK8C
Kpa6FvfVmIdSdLdKijxi4UJhDexjsWIV21zGkh4d9dCTm+2CutCvRBUQ3bcP5gZK
U7Nymal0cxTtfA/ET91O77FLnu92PSEdhJuwkCd1MnynwglHRbQ1SLUrjL3z2qw+
SVL+yKXrhgj1ixa9QHaQbtjzD0LimYipRJy8eJduTTI/SGjSrT+jXhek77uMAFCu
/nZjLFJwYMULsKFKnp3UuVOxoJIB6+Nuol04HuIap87lujQLPapMcd+Qrr1uv9EQ
bsPx9a8ogl72auQiyZd52LqIiKmfIYENqjG1pO4T5mvIMjn8SRa7OEk/e5bX8vQv
kW4BV3zmPCziPXiUf8Ny74yXw5a/nc+Q6ue6gRYGIL/cl4XBblsHoGZqPo30/bU9
L8ntrGBeGtm1tgaYZVp6sH6J43vYKYQoyxgSp6aZ3DpPdV4OJdG9KllsePvVNIKI
1WZYcfLRdJTveX2GDIFf6SsjcrCc9Mm/TwEu5tuKXcIZKRerQTegWJOXVqFN4yu4
yyNpT6xmBS6bFyhAFYi8jt6QK47MzguNcQOFFWQPfgbi2vs+TnzBQ4BoF5borrCg
Dl9xX/K3PFmh9BV087AHCF1vFiB9oW0r3lxftz1CL+sNOLG+mAsIQ3xHi2wx9TGM
zuNRkVM0RC5qbzV2IN+YWojO/2Gc7UuweZgt0RAGaGrwUd7vAQeDWOlmW2GcnTPo
dPFLXNB8q1m0pLCCUL9YkdXjhs9tLXFOgO7XSkIcgCe0LeistwMlQhBbnoJcUlM+
iL6F0BjuaDI87CkaUtMteqIFeZ4tnaGcjKjYUE8XApOPsWH3M3pFg5Zt/aWQPm2N
HAaOqif1hUYhMjT4ml7zKzdBMUXUcw3qjvwe7H6itCNNO/iNnR3YN8a3wqc6jb+/
kLLtoM/pbunWLUBTxqDq4hAqVTz3p7XrIch+H646JsmyJ8SiuSxnAYYEk9bUK3/Z
vVBQoDmXKQsv2a8rA569FWpq9b29Gsoq/iq8qgmumUcyh2Q0IRWlREinbcoJy9n7
gfYSdEpQoTQdbM/GKnYUWYsCr0/Xzel+GkUrQ9JvJ/+q4b3otmPh6CrmhD8n3zz8
mF/8DI1hqIE6Xj3daTP/N/yXCXj9MJJk8dmmcg7ao+dT1b0Jz+pFURhtZUi+yIMp
VF4lef0luh60EzaiZCqFx5aVJCPxIgUhtlFmq/qkOeD57APioP+ytxNHvU8ovfq2
iu7NT3FAwBLAInB1XytNnaLY1UI5CIJCO42yzMrBRiIb3MqpnYLsC0rGsaiqLkaw
CEUiREB0i1z7HLJ3zLn2IHMUpSGLk4Kea49W7xrG+oPGBjLeKoz2KHVboj0VWI7G
PAK6RaXiBvGad1zbU/bkXvhwiLfTt0QiuatNRuplPEvoJRDu6go19QYNu/DvfpV7
OllcULluk9ylCdPEN43zHmmWJsaU18vl3i+0fJ+O7tWtuyZvqzZA1kv7MiTMOKcc
ToWaq50zhWhdG0fkJqUQQmY4dBxVukdcGNQSc8jUphc8qlBLvswu8EcnUUXfHGiS
TTFQI90XfUs+wcTmuBTJf5FASUuu2FrfugFDs2wD9ZCsaTu9cMcPbnjh5hQIfaLl
MqHtvzPZlUXeHCO84N0hXMHn8NnM42Oybc1v3vi3qoTL53aDJ4p1HHBVRD3HAx6X
LCyOM0gUMnyHsXJDOsfpUWBFDwTqBGx9HUijC+baBVXYr051fVCEeGpZeKqB5B64
dENszgHdjID830kyiKpKWLV/NfqDDh1Re/hLjH6GxPeI/RB+GRd3feWrRBDA0trL
a38ySZ6mcCF8/Wwg1SS7CC3/2KS4NaVgRg+qnp5TlHxt4H1A2vzd6kFsKeVqt443
roTF35v68tcR89/Q+Ny8+j+Gd6Unvw/YOdf3yad7AYu1rn+A+opTlnTe6glHGDe1
wvCSIwF0gg4kw8xWb8kfhjmHCjWGV/rLqNOZ5hSuu9WjLlz+g4TEa7cXa6rHtJQm
trR7goCB1WW5O4TWdzV0ucuvIzY21VXqC5fozG2JSA5LJVbdiEnMU8B4pk7nOsL4
udgiLLfVESMn6j2g7a9+n+eBg7NWztk5dYydW35BEvKsHmSvmjVBKPo3XJ/DR0VR
dMTPzha3t3xD/ame5RINng2GgzkBMRoPxq9fRuihq6TBkvA18pxEb9H4gKhPXqhk
dJ4a6fqb6ljIvjX4P7uQKYTITXzD2zU9ihAM8GIA5K3FWKqyKQ+S8iFGXH1Xxrcy
dtzZjON0MMWd6TIyTgSw2ppReAjz89sSFuyHgq48N/KV+RRg3maV2GO4g/vRWIKY
XwAS6ZVLSKAVo3i/XDZDlFUnT3w0uXfLMCZHt+XTBT7zZDdiT/rvWDvz2kdnGAnC
LMp6GGdem5pnzcsJ/ahMHrvYvHuGuufB6YicpZ643ICJUJsonbpUKvlNm6Q+iy1T
SPRSWIWW3GwyuEXlFtjQq5q0x7zX2JwjjA4HxOtGaZON6tIwb+EbUFwg+0wJeoPH
pw49vwGevMgerOmmqCflTSGHVL5IIsjO0KGKv/swN6mQl3Er1c0Ij7bxVrj7niZi
0QFBK205MOM8bvTlmy90afBSeSxp+93VarSqzRDxdJhfWLasah4+xFoAc3SqrENf
yRC9MYe8tqCUhD1ev3fEiWZb+nQbg0V97RE0lHlO+ep/QKZc/zsaXlTNwVmVV/nS
g8G944jkB+r7YXaVWt6zma7qQCz12Tag2rSBsofcDwML/BxHImg9Rj7LfRQ21JDa
EhUh666XkI6BtfbojMJ0GMYRsMinfMg4c3vGUf1x2a4MJAwdmnh+o+Q2KvYEYbDu
6HLXv6le2qNuO97oFEpFNxRAV5Hl+7JIGzFTFyHBIm3Oe1A+9MdJpbCmbYcpH2o8
upmRbiN1O9SJB4TrsvTaN80A/SVHr7In0iLTye17swEZQHIYTbNGqwIKjo4vsU6m
2B4egHaEvsKE7SzcPrnPWiFLHEAw4eMy/oQFeBRpT1mmdTnLgVyWhymCBXNwKo5z
tYRQmf83dS2ZJBkELOXaIlxDyKf6bkpW4FyqRWUjdEKdUa8hwUEFmkEvMwte9de8
6J+0tqrU5jrONWUSaxQEJ7zBgjOw+KOg4kuPoxJzTYSWkus++QeX9nX/FstiTsbe
WDgpoywiMXMzN8wRcKMJmwks8vEKrp3XBKpuHnKJDSfpq1kxF1tiX65OCi2GRn6F
LmnQoPLNC1aSnOgz1nhlV7uQpF/2plry5TUp5Qu+iXsAufkUc90wGPOBZ35eLB7Y
JdYzxeVh+Zo/FAK6rLGaldcP65YkHX05xk7cgRbE0By5TAzQ+PwrMkz2LK1XFYvm
tP+mlxfrlfymazffHlrvLAfgyMqvEzeHDCovBPUpVNutk34T0H/1g6m3hDn5JTv1
SW4oqLIhW+xTHdaF//j0IQuoQfFfHhyPq0WT/2s7xkPHqzxOClDx88J7xwuP8NDG
vNUt0UW0/IAITMoNtgFVNbd98tiWjf5D6U95mnBvIq5pQwXcIvpt6fdsLiY/3JzH
Hke82NnUSg1uPlflor1pM3G3kZffJiZJlSwDouHfVCa5qGjAIP6XP3qmNC/LHYL7
SZS7IdbW4ERzwyOPzI9DDQiKS3xCoQqjre/w+oFnjB3WVnPDYqP/63V2Ry4+tGlW
wqMFyTIm4xcXGVKjj4yctJZQPRT4RS1tyTBKTnl8H3Oha6Vkw0HozZVSxW2n/EFC
PDS1cIEJmHJj9AOL6Owfst1J3v7DUZgXDwCKds1Xj9U+fgX6rHkICJqeDhTXyhsg
/HJshi5FoFZplolk7GO9AUMNHI3YaGYGRRtC8qultQkmMYfNnOJlrBUwo5E175n7
MmLsvW4K4AlawBw1gVuSETX+0JapqCMuuJPKp6b970Owtao9oKSPHvRB8qei+g7T
pNqujFol6dmA/91GVW/lW7ZDIfHtMq69VIhu+3QWFUoGItie0ArZgenrPCr3Tqfu
tvXEw9Kwvty5PSr9H8MB4P0ZlFRXYcb8UTQPjXLeao/qVxzvavsv7JstvGc2m0FZ
zOJxPv2uuz9BLRaUlpHRVEAurIcmv19ABQtmFmjmRZLIshHHNedsHj7H1EBDS3l3
3JKLNrZ2SBmG2wSBpv17wv6KyOtUsT63eUnc78pbbt0DbIKtwXKqce4hxjYUoyJT
oGfk1EGt/WrVG5KWV7QI/w2Qw98cg32UwyuHzfB5vrkNfj9oPEwnGEIkyT6OXGEd
UD275sBjIF8xOHUjVbAwYt+gvRXDsFnKYrS0RqZgzykLkFV/drbL4r2gBrHlOW7f
bCwYBJ1/ZJUGRBWVkhk885Fv0T49d2P7ZMf4BO7jr9AJR/16N75LSmDvowJx6VH9
k3crZxgU5q3ouDY5gBWz13LJhqPgSIWiZO07tUXK452XV/tpA2MSQzbaVCyYOHV9
/kL9sG1eOjidR27Qg/0gc1RIfxTWKdiAi2Aa0epcdiRdvnxEpWbePoeBq4iXhGGZ
dokvCbyhsODEvda4TWQp44ZKplS8947sbdliZ0Ld8aZ9nlZd2rnymIQnZA960z/x
Qundfjhphmacq5dKyvkFBmsZHp3+BMuRrhEj/4g9U1h3WVReM92FQ6V2utv1a9xS
LiDFkeGKq8P3msHQiQppYjIn1Rsdu73n1YyO/7kO9490PDJkLM/4r3Sx9+eCA0S8
dsBwt4ZVOxxOwvLNHdIwQ5Jh73/YYeZ+V9Rlj1fCvX1CTAw/3GMe/gCpvr73uXT2
zC4oyHKlYdbmzIreS1Qm6NFUVWn1iwrYxoLrssxn+nahkjbQ1UIH+Oxvyi9q1jel
GGj6MF3B3ugEhtBph9l/fEr53E5sG4m06QhUGIf1geumkBd2aqMci4IeqeTy735j
+nFb+er5tYpxyUolPfbVUgnHvOun3a2I8+GoLXNt4PIsPuyxF0hN2wFvRCrjAU00
tvnGV9jpcj6S80Qtl3c24KwXf6BxvfrQEjRx3Y2UiX34/SqssbCPL0gDxb1j2Ggl
sKiNNVSiqCd7vgi+0+CM1q8ax3LWb9KgKNj+dH1OczSSGGtRe/9z4jkjBnqQJfOY
PMBFv/WnjPmlZ2+7lSKeXIVh/SADk/lAA5siZM5NSZmuP0JzpivODgXF8lf5TW7m
SWLCyxHm9L83j4ggGLYz1OYVMTNkVVLsG13hYlUTQEV3XWp8ZEqhIV9YBPzi6MM8
n5hmIXIanOVdsG0QoBG/+evHYgt7DLyILGLXlF9up0qHViiIGg+7z85Y87iB3s3M
qb0r2wTye2l/vncuxaeQbJgEf+6tSqxc37MmZeQSsM89tBeyL0/d/rIc1wtzXsOQ
3zUH+dIB2q6TDMDlHpCUXqBrjKHiuSUpLJlUJeQVQVB4glmHbEcdgkXNeqvRaH2z
lMJXdArXqyj37UTQXhvAGvied6WLb7fV6FWqEDN/hhpGHPtkWu3UZP4m5Ix25Vhb
Hh8xnqqik9WzhaOJtyR4B91fYVQtT0QwMHasp0CiNdllXMcegJD/Bvtx1SR+r/DH
3QTHnFfsMFn36W0rFAiCbZdgcqbwwqDXzy2jmdKUjuuDKe11cY8Aq8gVhUhQpGp4
V9w1LCKfVMD/XSx+WLKaDhS8UXOY1ns1ceoMkUZHjzBW+2Ty+HezEvUI8j/SHDZA
qZfO4JcwhbJQ2/swGhSjJTpc3PVqE0CTnmtSYSnQt340RhVe+K9SQJ3jVOEwr2NK
/o745cqNhBrdH2OeklmjgtfzjrA5+MZG3HgIxfeKofb1Guo59HlXpEW1Anw66CE1
Ij3hdyn92DvtZYknp78Phme1uKcJEtAURHy6Meljtt5YQayCx/Rps8HUJNLFY78E
oSMYRPclN7zBy4VPfRDZGaKIKPyaNLJeTD/OSnE42QgiIcWyBgkU5GgN8gSnUC7G
HRt4btPg2g6eyDKzlYkehZf1+lAby6i4BegwjcJUuVuptGIycJiQ555amgogxe1T
rEdaJPsdvWa0oRV85QBwsu4mJSgzxZwx8yKTiLBzbcnkq96TAsilEXkojP525dAv
a2PuM8Ce239OrI98fxJf0xDT3B8FoiTfHZ4RfrowZGkXFYN36Cje/jLh/daHRo0a
my0+2PC7PEz95nkq9R/wbjD1nHLPXRnKDm2fXIziAArbcR6/LaL0gyy3b3HyHR5s
gak2jA7KfCMt8rGR2q36z3ewEUyiPNRmClA5yiVLBEdxmxRVEbYAw8rmd0hSBljm
NdFvij6y9V4bnll4MWPqM7bLhBAKHFokh/MB3gRphmXioebBl61xoE6zX69lxfHH
/QvaeUcH2pcvn3VnzlfHR5qu15KW9Bc/82cN4LT6GzvnaStjsYt+Q2xiFtKQrvRB
BG/Lm1VvouIvt6L42p2aAyqrxq+cyFvMHnH2DQKLL+ngfKi9twoW5QsQLeTV1H4e
4l0Uk9LKn61++rfdIleenqBND1FeZHmNG039LX+5eBAFn6+c3+hKTmtQfT2a5y5c
Qv79W1Ey7JIgwJUT5iDOi5ms3azHgxU3lHhSdUi5IPa7H60XcUSIEo0MXTOweX6D
qcauDcWXuPnebSZBFny0leWoU5E4kNTQ3qKdroMzeYc7I09SrF7cd6ngg665ltBc
Y8+L+gEKGaSVAKK6/vS6GiXdrQ01CIuByEOh0a8qcZnqxAI1ipWI3Dcy735UKb/k
ROVBAqoM2lF1PpsVE0vQmNsfbHaxkqKjeS+vcsWC6YT2GtFFSCB7g811cy8e2Qub
3hoNpZs0gKhUgLCeVF7Jxf2HthJ01WqhH4X1XtEiyKOepXVl6U9Ng2VQ+gHH4sw6
fYXvGcaFG0ydc9WGw/bvCYf8ZIxjFRuEUWOLxDqB3x6HEHIh40cZpqYz8xeNh1Qf
FXr/yaI8PnAVtgF3JmiI5OaalGc6rgkk2MoseGlwxZCKq3wu+w7HzdkAPL+vfzN4
wz4+s6cUNaxt0DdRzW7sZQMeWRxTRQUnbn3oSEokhZ9fbNc9Tr3EA5tE0M2LmB74
jLTdIAA6KEwHdZBbGH6Exe63lCB4e894P0dDFxrVXzb49yQNm8j9mASLcUikM4ZF
NN3MV0oeOZjrAASh6Qeb2yS3WGPQJCuYFpUcT3hBFUZiAvq1Q/GOprn+kdSOX9O1
pLAXb+AoRn3D7kraMR7Myy5+S37WlSa7P3XFyrlr0zQnNw9WBYvYMljPvyrMi819
332JNIGpNIp79enDLHHlwoHqgbZuUJE8mdWAoUTqLfSz9X3HRZoUVyDHjWeH9uUq
cshDxq3/0j3aTEHdM4kf+idUUyPEzoY23Wp2znKkiRc08JER+iL66/+WNqOLI3ll
A4znzevOsPULCOuLyuuSbq9bgk9nTYeDxaapCjUJeNERHb39sm2gaeWVLqb6b7/Y
VhmYv1fWZ6XmCBqVHQd7jvKWULyzG7htqEsA0kAOZ5K6se2dafAHrZSVTGRm/yZ1
C9F4Sr0R1zh67Qj6bPemZHK/Sh2YTv6ZircLqbssoca1GH4vZLASvoM9VmmVzsoO
D1oDQ/MXe/jzRt2pK111637o9byoHIzCLUR7cx2kta4hX3qCSS/YVetc49tgEuhh
LYkXr7mbmbLLl/zFkQqdwOiU5nUbndIzrR0eEa40bu4T9oTsEtHhTDQuseARTAze
ryRL+siUETKLgV1znW1eV0zmi6Fbgrk3KQ3PN8Ckim6yHjwxm0TE9aiTafJ50R29
AhFwA/HwF2bpgUM10tfvfVFn8kTB0I0BGqgxroxZ13kdXGIHF0q90NFcYWC3a4fw
ErCJvc1BEPp1Dgr1B3DRVZ+OXrMpzDqxJE46HW8j9ucnDTvwStsri+yMDsoOkh9T
cuuTkf2AgbUSVJKyZgotZpHtnKTWBYS6J6O2CTFRYooYuhTmlAP/R2wlpJ5Bi+kH
bgjHlcheGAY+DdDNThXyIZKYh2l83Kc7L4LTHu2RvGqR29LgdtyPezWR39RwyiJX
yNpfN/a2RY6T+L7arERTGY5NVSmoeU+1aZ2KGvBlNtGrYShlzpWO4DG/R4ev0ChK
/hrRVXDK4VQuoARhQxZIY8WBDS/uDUx7E10gVMuJQnoyxc8Zv31RABkoaFLtjBt1
O+UyVHyTzKb3dxlyZjiCVxf0vgrN1zk0S+FoUcCuIfsG/XQ9SRyaN/qCfzRpze2d
r2Ir0z6/SzJbSZE2rGH+TCZ1u9KJz5edOAQmfipIxGPnHSe3Mz3jYPCUKCFBExYr
j1Q6QgDURqnMWcM6lsKXkhyXeTRSoiouB/QEkzSXdjHE5ZVd3b+bw+Om5HuO0CFT
aONXg0uIJDZoc3Iuf2lf6kszO3X3hUwEEpgSEnKN+x2kAyrTkDqFPTagSqPnIv/V
5G7D9KNEp9Ap3I1UemWuAgm98ZosDV+putXmnUa16DGHwbKTCk6NdsODLi9jNDlt
RPQmiACsrHQ5EzAwXdZVEj9W2x7VszKqVYpVkxjyr3IqXW4HjhS+0yI3ZxYzsHM2
pitSHGFETYEZSAGM1ZQ1MWGwHB8lqybSbP1lSHjOY23HMSJSBhTNhI/T/s7mA1n8
AK5QTj3/4KvoPAsYEfypOkX3UhlXHJLMoBA32iDS8jsJ/4iRH8CKtbipHNPLIo0U
RTeiRBYHCgDZ/P8gLmlcb936wnW5YUysxcGcGgfXS7Hk93K1qm83k1LmlL2UN4Im
/D2TiAgVpZSaqdYxRgZxT4JyUnVlGoRg+/FoHtaY/KjocCVTYNQJCqwUqCEJaUn4
gp3YDmIy8BB4N8ZbPOK5ZeNqxSrfjI1SFKFVIcENuLjipvuIQGlYSipQ2ndvyRJi
imPPzpQHqxOIsBkim3qf6iQegb2B//Pc5RY8gHdMwZTBXC/r6YTlhe6/aZdeHOsI
nhkDToUrtjMz0gfvZ0EWV4zH7j6Z0oI5UZ6EpctRsroe/btWiXuj/n1XpTEAFyZ/
S4+CQW+KO3qDuc79fbUDQ1Yp6KFIgVG+UF22nqwpZElMl/o/L3fauf124qOZpIIW
qo2te3k2A4tubQhf0r0H4l7WgNGxmg4ewABGpopxXYsit9csr5YaW+xo3fR1hEZ2
IGsbmRbu3bshb2FMFgJD3swknqxSjVze6U3gnua4Ji/IPWwjrqXaj5AxlO2zsjrd
Qadxfo15BrlGKQNPE4reuMlAGiPAO5//+9FUWsm+4w50eNy1coS6FSUZgjuLdE9t
XU63/GG3y011T7kBLsvRd2SQUGGgzd89ZhnXCnGLyj9krWFZ4cHmT2d+wm/aM1Pb
f6MLO2noEK08HRUaJdFrsG8+wstJL8hIuu4m3aiDODuAOCJdZhT6/bknvjQ/pqI2
LWqpPDlkt4CbIhDpnXPTEByqMeonLSk1hvXBBgOUBR9OjFVEXHeC51CJhWN1Kl5q
iaS0EQi273NKIV7o7BKOT/oGiS/YrTZG8CFN7zQRFZOKM+qaQ4jjLg3vWJcyPaLu
DY2PFV+exwRd6imrvjsjANFQOE0W8a2i2CioXKTl7lt+xf193/+SVnmVFvJaahMZ
tNkSKJpsiUkEHKAadkrv5jCkpGLmLlQ2II5G5viU5iCA4ENSLoFbX8sQ0Nk8qBJ5
qrUaqrUa64vLQQKjzXQvtZe6yoZxOnrNFF429DhO6NAjExpiyQm2UX6lwnzUDQqX
70+sH81xPc6iRSh/60CRbwu6PZYQ/7lCpENZEamS8UuDfh5a2PLH8Z5C+gE+UeiO
QEf3GYq/uYRyayw/ORDp5hUacSrdFAIL3LgT2fimd6cczsyaw2VGUYeybwiFbhi/
VvQSJy5Mwz7AFL7OkM2TrdFCDA4jAtxgk/Mm2qc65EoeJXeN49lAudOeWHHdKnRM
Oe9Baap00dsD1DnI4iHDxQWrLIiKNC4MuSOsJ0bW0lqWvKA30do8PGEtsQNB+TMC
aYqPTX9jhuxkjyCqlnjVXT7qlHymLIHTeQqqOjIVa5d+ewCK5Yp2ttUKHhfHVO24
DtV2QJFIJVuVpphq9jkFc5Pvz7ZS6an6jkF6l4btxmuMdiRXky33uaHOGEi5pd2L
pXHnBOZJAbdWQCd25/yXCfVsbVcHa1P5iww2i4eptVOXTohnvzS6rN8LbFdJEws3
WcLKDGEISDt5tL+By1uzUmgN+4FVc6EJQ8T5yOSGXJZqIKB3azhurd7Z6OZ62DIE
7mK64eN0RToD6Xvv7qQ9+RclvKpKFhgs8Zbd7Uo9ghvMlQASKqCRcdqvvBC/lpeH
7ufOidyINq4aKQIuLTM1RG9cpjqnLFJmGiCDlVCX8HCP9bZGowqx14A9Z8hfDl58
jAcg3WwwmgGQXNLlJqJD55pAFNTUWD60hijZB9tDw8KxYhTkQtDsRVVC7Sv3cJ7A
nyYOgNaf6K88fPQvq9S9x7Kqumrh+BDprj6ZM1dnRG5k0mf/D83q9WuxWhcJlB5f
JY/ETV9RJIlNg6GgFbTNu7CE9USjySBb1NBtxlYgDpF3QG1TEj9j8espQ8ehEhkX
1Dp32lWTFGi7elG6dvBluDa7zOZn0UU2edkMPQHBULUibDK2gC/mU4mXAkUhp9Og
Vc9DUYF0MRV2VFOSaZJzbguZcDCj16DhF3j43ezhRg/GfxgKvpS0frqTke9flAVL
N2uMN6NmurarecOG6LIcbxmQp1ovY3g1ReUx4TyW/Rh8dQ6oJpZN1vJRUVL0IGKh
TPxjHa/XibVHa9frN8XsRle7KQLzYoV5191wfJ4Z081Oc9FwB/T50a7lavmkUtkl
NgMtoPIPoTl8misI+dha/4I2N5my6mh3NwJfd7fAwaNP6/qRqbOV2VSzfz8rKrl9
H22p+Rmyj7nRlzkI7E0eh2IqhOBc1/HXlGrE4e0hyIJSdZ744ioMlLjXVgrqb7bh
iYT7AyBHVTS+TTYpHEUrZCiKppaTlQ081a1/3kPcc93dihmlG74FhfYM3wMVX0pg
y3t2Da6QOslfRny1DkK3WlNTg9seHYzMioSbYu7Ihv8S3PR5FBO67G79ztlCwgh9
E3yfJWuKRxWLgkZlAhYpaLJQbCoO/eQrRcAHsUDXDGG83oUnjM1IypCLpl5n2WPu
+CNm1kLKoE3E6MyX3aXwEDKRq2h80nbeySet0awbbvFMU4Oa4L6XRrezg8raFcXB
JWThShKFGfScuTHC6gosO7SFoFccxs+DD5VTI03sWvCH3AEzVo189nCBKO+6mPOA
TrvN+IqmOUf9CmbnFXN/MLNoTQgAvH/Qp+1pJIKgFDyA0AWxrCl4EB7H83kGS9qR
MJKZpoKzsINKj2eeyggE/9ILwnG8PiMHnTtA2Fras+/Ca0bNPsew/obtaA0rE5u1
HbK2v2lxf1W2cuV4yoRGrVvOEtfs8Uc16crgafRo8SMFRnh4icUwkzuGei9FXSHl
q+ciYO32oJZv4yOcWel2M1vheMgLQrdGTJ7ZeCeGdxr8Emtab7eRXAYn+a+VBzND
EYDvEEsXvZNwDwII6LZzrnTazD8UbMLWQSu3gvuiuT05KRl7qOsRIia7S57yFN9H
qv0HkdTbEBOBu5g2ZEW0PgNZ7crXDtjXtJWJ2PetNpkowTyCqcihiynyWcF1Tj5z
yoQQOnsSkYTCX9FnBVzxRphO+NY/kaxzp0Sor/tH7sdGq3a51XvBRH6C3EWP+zNS
3ppycgkYTWCeykI7Gnc4Wr6k7Mkm/BT6GcptF/Zyy23q5A8J5aNZ3bgvWVwkC6pe
5pj9Jv0+4XyZzmHjPIiqLSxFhgZqE1Il7YKkiQXKGaFHrJe8KCpNLOmgMBr37XQk
6OInGziEDOKRf7I472Jj/dIJsIb0FiABTxymaD1wWjW5Te9p30OBPurReKrO7uaL
WifJa3lHBTpY84gKySxL+Bc+w0BakPyRSXQU77TjlLMFn1rm2d+4bRUMHqcrOE5m
ctK4Q9eD36cTUx4j+/u9/8Z5csb+UEqSJQsLFB+di1vt05SWRcZ/d42OWM9zHq7E
uV/AEDoNdBNH+g1Qmmwx3AvCSpbZ58qA7pRb8w/81M3Wm31My4uBgk1vh2Lak3yH
9uV7SAvOfItmKIUo9wcstfX8AGImETiijcCkr1rTj94WGR6bBWzEEBFtutcckeev
GklHxa6ONihU2NhuohdI0JvQAt9Atz1QUCtIYeMRxotW5PHRNUUev5d7hhAm9dtc
Q9JDwqG48Q2FogK4XwlYMdQ5p3CYIJeDFGYn6p6wqVDBddwEyX3zBVcuC9zRzJVQ
Yt5aK8icaXF8jisO2lD3mmywN+lBkLoyfJ1jpK8t1pXatbj8NpxwlDLpT7o9dBdW
nnjw+ZZt/R71nqgTMZfbCcG4wm8OXROptf+PYZNa/E6Ms4i9sXjjG3o4zmhDna4M
weX51aF09g/f4Z3x5iOHfnGPuhAg+rsuPikf/031RNsx2+7PV6dDLTQwXHrKlFWh
c0V/5Zo7e6etEOVCgyAxokc0k1Rnta3/2R8iosDJrakhaxLPcJmTWXf6TOEi0L2C
SH14CBvyjfvmV0pjLA7uU/RgmbgPebvqlZgGBhHUgE99JzGxRwRyhUHi4fbpDx/+
WS3wNt6lk+aNr/nxsxkDBv+fb9/P5Tk+m9Pmg+LpjVrXJRVl1cHWw7YKQMWNAiLK
Bx04dPqoJZA4WTnwxxRJKSGuAHpYoEL5jim/ccuINp+PkS1LWc2tASE9uRWlncvp
fQeVKRdfvgX1tidyBeLaWUmyY2KAJx2Ix5AcAzQxbP/VOevIifk6+aPOIFcaBnP/
kzRkY+bsMOsdG3qe6RIovoO29jfrxfFGbI+lM3e5VRFY7KqxU3RbWrQ552ml8Qfq
o+3EvolfLC6xTqKfXvS6fh7MrIAQrY1swOcbgIYULYAuG9oaugzlV3erJUWpAP4M
S6IdsvHdFXUhgBC0b619soePQWax2MYIkhOkvA92TAKStsKEFQfFiNzJIgOIs7d7
D6szHdXYNMCd48HubLe20/VrV2koXsPUwwNT25BuPWcTUp3+KOY4eIO5Y6j4/5vX
02NkVlQRqK0W90yILWd+vVFnjhPBVYxshNKmB32CLdUI8GRfHA0ZUDP8Ly3wy5bW
fTmeBDoOEGylbvYOArkSXNFFzCSUREiC5YCfHWiG9ImbzxNCDcFxIBj32l4jt6CJ
VWpvklHyrhXegO/6z8wEPeD87JaoZ4oqZUh1vzNeOJR65e8Pvv4GJIECjsx7YNIs
9NZusOwRcL8i4QyGcY95paeyplVAAUUQnGj2r7hgqpyic0CW/lHEeQ3hjUtnlLDc
EpVdc5jMnUhk7aEhVNBnqQxiXjXSae5RiHljdKPXbwDD9XQ0IY3M774XF6a3vViJ
n5q5D6KghejRWU/NRFRTkkh0pNwYtkAWDtmJH/vTI+HBHcVcFHs6TJR52D+UEJwP
xuQ79xsYyugWUCwEXcQL8+aIoaq9wuD+t+bwm9aXdS5RvggB/RlcL2yL8eRZ1mH2
saG9ufBYtnGYvhZfNnWK4bu8juIKTF6ctOZv5fmujLXOe91yZf2fYc9DBdaqw1zx
NZhFSpHN6Xco0t9ofizr9hP3UcMHVN0n9lTuXS9vkz8sX84OKnALFmsv4Eg1nzR9
I4YQ6nvsMv6RJ4+xFKrGOpczeF8q8OzqHxMlLvnu3X8oKNB5Lz5+SvmQbgaHPipH
hhLW8/a/VY1DhGydk0w0Ilde7dKAsKa1JrTd7c9jQZ04lGSZ8mScO9fEaP4cx1Zq
yBMgzbdTS8rnigrNoXfNdA7hba0Drrgu+Uy4DGv+GwQosX7rsLbtnTKLsdNvN+YT
S2PkSRB47ZfkZrn+vZ5OQqbRAROgRMFuZ+W0f/jZ91BAnzjDufV73uuNOw9NPVE3
ovOjHMnz59euKRwtZ7xVD0LUyABlIYNmMh0W2Q/4L3uBEqqYEKe3FVFvA0whNJtG
wFPZdUaVsQMD8arNDB7aktBfIQ+PpQRhvQ5v6br8J51FEandiukQu+U0+qT/WJEn
yuYIFGwObTBFSfpgsktad8ZQaSjMNUtRotDg8g5Qd95vGH+6fZIj4F0uvLt164l0
QcT2bmLBLqkkfI+nonQSBA8w8UmujF+pIUSGTnxxkSq/q/Yc+ABEiybeTz662Cix
dCBWqj9HRftZkEhYFrI1KIwgltoC8aQpue8PT35eJqHPIYVZiDtxE9Nv21pExOFT
3srsi93N06yQ4u3cvVPDkMIraiZ0haB/rIiovph9kVwO9LTRfhbfQL1uCIajvqJr
ifEJyRKLw76ASBLKOEAVknU3kY4o8jzXEnNONwqT72cHvJDiMgHhU1lxNsBvHTzq
n1niwfcNH83bIkfnuoAE4IUgMN+cpT3MmUJ99yPsjXAuuOsGXnUJv4gCbL2J4/Nt
I6TX08fKsoJmWClT6c/PnMaQj3qegm4aEv0cEy8MIxD3wMFw3dxv6CARcBRXYW+q
27G8ByLJx3tp5Nfip9s68poVG/wWtkNq/T+g7xkV11CEVfMP3nPvup5RRJsnBHBl
DUG1ohKK3FdEIVTktdPJ+KwcbycuoTEragJbJpJSL9pmF5D11TcbFiqFty+3Yhnx
WWUJn9iPRO4xDZNy0wyAUlU5sQL8FFDC38RwDrncVB5muncjh7ytIbXM/r+Gia5T
FQP+S1I1AoOnr8jGea+0Rw6pEoqLlO2rR4E2EEr9ioj3ev7k5zuzPaFHj0ixJ/3T
vGxGySzb/MmXeHCjml2ngkwTpadUTvxG3L0QAz9LqiIkn63F1pfvPUNR4uhUhHnw
c3Ky5vcm4GCSmYi9edm3Wg/rK8KHvY6z9wwRXzOD4d3pfOCFY2K184ghyzhxr1Pj
xNIuRmZVjHh2PeHDjxTM6tNgNdgmqlXVAbtffW8Af+whFFiIahhE5lnp85oJ+DGX
iThhf13FA7A+IxpXTXBujXWPijJ0bmoml0PeN70Kbiv2k1ocuIR92YQdLa1IgygT
nxE5D8Du5VDSRCGf8I+35xh4JvHNyydRnerUjxHxaRJ3txO19JrbxyRb/1otG5eA
kQWWZQDgga49p9AJq/9CZQufjuush/sj9oyUqMdlWUCGqLIsOI/VFMyWRC2B196s
qox8HRVOxuz2piDf6uo05v5X8EaYKysJCiMn/824+fi2WzLie2TfL3UEuHyyopGB
t0tDRElIyPV2g2lEabi6C2/GLodZf1amzH1NJEfS52QSwvirq7VYCYRvwi7djzeM
VQHOseyOqfNz/XoW9wA7Ydc0pZp+D6JKPCNamPpntuEAyvwGvQMoul0EMTlY/sNS
N79nO0EfbP56Otph3axXVTCpdt0Uy9D4+5dXVdwLI9wNQvMFknD6J7HjL845vQRx
oeVzL43ASwpgX7PK0gccA0m+qa8gQWOEMowoG4imNTmmLkJ4Kp+ush7FT5xrAPGZ
YHvcNbJ/hoPoplK4xYJ0IIotdQDiCJhmU3+dXDKJAMI09gGkOnfSp2870WwEv5EG
JOZnsGVKZpZERZjhL5BAeBUZJGaYz2ddubsU0COIgLJTqN64Eyq8lPTDJkEQrEZ0
yxMKbajMz/rqczRnE7BlIuKpq3e7MAh2hXiSE4hQGf3gW13NJ8tYKhJpUDtsgbAj
3PZbUatKoF2ZvZGtLrGwkvx1uIhWKUaG5S/zkfGaQH6dr8NwejQKJTWsHi0c6+u8
i9smcR4iTUzgf3S5xV5eSmeYrR/XQF/p3Fiz55DhabLsM2KhnhRj283Jf3qWZyiG
rj7uQrapuylp3Ud9EItHDy2AdRznl63pb4Wgi0jAh0V5L9iGA3Dzr/QCIRMuQ9vl
bhSF8YEpYnRR5qz0WZkMDvXnP5VtXH7BHnQ1rEzweBr5wGjPbxS6vOkm4DUFk8/e
7J4UwjxQ3Nprgzi7RpUUvrESx6ucpFFNjZhdRKJ7h3nIFGi+adMf7t1HrH4QEYVI
h8Rg1KxsK4e5i4Bwf947I0psXXvVnOCkV6idY+g1Wa5F9dtYYOUcR6Ih7axlBL4o
lVXUksm2bJ9k2eEuvdB67PSpyi0UWyhGm4OSYkJh82HhSU4yOyHSkHUuYd11pUa8
FrOzgQwV0YccneSQ6VPZnetlVTRJG8EreaMrEdcoeOah8nqmd7wbFQhE1jgvo1i9
yFHKSA4gcO7zSD6eqHutcPPGvOHIaMovZ2MnHvstfuNrYv02Etvr1XsXeHde1p7n
S2G5iYlCWSPD+vUVcRwHZ+Fpw/isr6YeJ7YbDSHDx+ttReyHdeIL/zZb8yTIA5Oy
UYFlTFxUCeiQtMowF1BnHyxqsAMNDdAFzTXUreIJCZW6ncZnFyBZ0ZwPvPHpbcqC
atyHt/qCc8mJ4xqrOvtyowc8wD4yCS7T3+1DKVnMMc5YMHPd0LwqYO3lCkbN+IK4
pWpjEj3myuH3DHfd3miQw3kLQM4svBjOJQtC0mX+kMdPV3fyEI8EtnBozxd7rsQF
lXe6+3ThcH7iYISsUd5aIzci2zOdoQgj8MQv1+h124gMCF77TnSppfgkrHAgqQW3
3ygUJ/Lsgp+5oHoTpYmO7eoMY5CERpb4edYcqMcoaJHp7wtvHYYOh7UeqOZr0MjX
3+V9rIhOVANo3FFxe9ZC2PkYFb70fSBW9H02LyMxaDAW2kBYKeAmDE0CXWVBhRuU
71zo8mAGE/USt3s62KLGuLNWZCpi/WfKdw9YsC4uLpCCg5Bb3QvhL8KtCQLWy7u+
QQ29OhNqjwa0Ez+LUltQE2DfpHOJlvWplVqj9rRnIOgK0sJbmL/RkkptyRLvKbVI
slGzFR8IvU0i4DvEPJBB1o5ljg/A728vzzXIgyS8aK2+fmRzprtFdSWg8M8Ppt6X
SK1dw7btKfJZcHR9z0xp21s8s1Y78A9zwqf3DwLhaZjolInq5txbM5oWeRyAyVZY
ItEheksHKVcpIplu4Q0l/vECvhGBu9KgKw8IlK/CCE4AJ0NSor9HxAhg1OGL4LZd
C9VpyxlzrIx0ANyCc/5pvnUoxUE3ln6sFVP3MTgjlTMH2Fd/XF0f8GksRdcH4RCS
wg8rh2me3YyJc9zoc+NqxE0hOgeYE+qEu9SnlusdnNzEqWoqt0AZrAerO5T1bdcS
zilGYodjRKln+p0h9n7IaZO7MvS5yzjmkdKl8YBus8rbW0YQKk9T4rGDAoxjDh/E
R7co407tZMZQa/8OEGMyo8btBs5G4hLGPnoUQ0TGvQOM27aCy7NJUjsGdqn9te6y
K++72BWG9x97CxHRLZ+iR5e5wTNo04Q+hr873Kvmya3XoDQQHM5QJbr1TqxF58cY
edTMJErBOoB7Rz5GbP7akIszRkJ96TQCe4+nTvuvy0iezH1cogMEWPpKj7VNmi/U
aYeESIqmPIah39qjkebxOw1ynXT8xbDqCMMOO+q1BjEHiIhQFeTHD+YZ7MQzy5dC
9QrfWatnqfz/5ovQXkC1M3i0Q2IpPEl5w8zIpWHSAd8Py2qOcgfdu8RdCz98Adze
AU2MGglTJbkTtkFtujRk1xlqPlgYLJEzwaQmYzPHM7lSxOS9x3+kTmtz/n8wxaC4
68LuQf+l7VtB/PyQ5s3D4S2DJqBu70+FmZwhpKiZ2Yg5ISe0uAsKt0ThcLkTQs55
Mz61b/bOxHFuGuoJzgsyk8lWlpjQrPhl7nXbxqsCyXz3FdJQ0eEf5hHvNuf9gQTx
OeXGvAHpgADjq+r9Tq9abyd3ou1SF9VK/5cTkniOHTZRsw9wLCNyVlhVW9/FlZgA
oFpOQD5UzV4RioB0f1SLU3c9nl8pbEk0SSJE3sR6UOTO0fp7sKZIzr/5SbmKyIDN
rPHXPh9VvujblSxhmSiUgST4YdHcVgnYhpBYdOtVCxryI7RAWAcPS5wsAgYiu2GH
wXolIIPIrIgYLqxJWQBx+LXWh17fiABvxTKXPWWrLaKFU4Jr5mUnUa96JTGjn/Ga
+VaJ5/Sl/nNznAg6V+tuwY+45f+d1PWczFLU1gtKmCrlobpkcjY6iLjC+VYviHdf
FZvyndAY6tPJn8tBablA3moCLj4yRbURII6vC5r8OlvrURwzzwGoB17b5llpgLif
QkKykLtfwiQdH0Zr7PfzJtBnatulu1s0srdHH/p2Fjk+Uih5Iqq/RXkGQJu6FUBq
RDlEnqkcY9g4dkSwtcuM5E/t9CcGmU3MJfUAsD8xT6eDTbsnF4SrVWX0mm2+MSq1
CvIfILiwU+sWDiK1zIWY87TD1M8UJCDZMcQm8qxfJH081otznxbCu4MiRsxp0L2Z
GAwU1LeZ2LD941tBZF2lKpwjcdU91+Wly2o2JwB3MJ5cweJtSewj0UR9ZBiiEMUQ
peQyhl8O0IsviciVOyOcrZC2yCz/ni9LYarT40JTr8IfWhXSYv3wewzw7swImTRd
JbjelcBQQQ+2QooSs9wTRX/dBqzKK1P+Fvb9cAV/gqGu5Map7xt+1dv5mrLUKq+w
niGTPd2gMQhmkhM0cMsiGmbAO4uqImp3CpVMQWVtXS2VfY6ozIDedfo2GzhV3j09
S9FqxtPxciNkO4ncngf6UFjzKQ0DBEqiYzT4NiiQEIkmS/BXviwotrNxC2iBdaeL
mEFaGN86ZlNqemiNKYQXLykwz6tDQ3lzH6LY1iHfZvUZ9kT3iSniURSj2fuiFtpB
XrtC9uf8y9v3tzzuPqiAIssM2rjog7qUzEF90Vte8uILWSy4+oIWJN2jRRGao90p
622TZwLGX/OG8597kQ37LhGnleHKhokLapmeNsiYPh3UFb2jA/TWS/JtyTAZ+c6O
PwroxI1y7gGrFi7pa72NduCfK0BRn6dLrhbUQvzRNal/7o4SalrFhXpLGzNU1jjb
xLX3r1PCJjJxzA8rK+501piu4KRR4Nz0trZFhpvKfp0Shw1eY9nSTUbB4A6Hhlav
+KKjwlxBftBdYWyj8/8GfV6cbbGX1Tri/2YiCVnTNF5UySn+IpMLncBSZxCUf8Xm
o8VIFbWC5qgwofCI7PSh3tU/Sljvcu3IMgxJwpkRE7KiGzZjc9+B8Lh22DHD5bf/
YvbNBPPr1Qzp26EdO1arQ69Qkni++E3XSVYk3ZzHTTDaXU1VZcMRS/cIvxERpiiT
N3CnPHOLjij4r8ltxnFTEmQWSfSF1W5K5lxJJwb23/hnQvpmZDdGEFTqLGBu0W2u
HryjM1zVPsNa18SjzV3cuw4GWD5WeQSzDuuYstg6ZW4bTKpZnbOBiRfM0SNnAvMo
aV4gRsof2pYBHE9qA1/GMbg426F7qhOAc9YU1B8qIt12LkbbJuX/pLZD7FxyLEDF
yTV6qvNFJwyogpM92ndxTKu5d3+pM6QQ8lSVxLTfcwR8sh5fOdfAwMDbfLyheYzv
78PTGyiqEcnAn/SGg+AwyIlwc8JQ9t3+CCLiWWAyv2Cq06QHyB7FrzeKfBcXyo37
vtbcNO7pzzosntcHzy17DT+BKdtFTK3k0YkANAyyhOHP8nANBGtObrfreECjuMs3
9NKnCCNxVREMDRIAQBnlNnzWb2gdJpLH8bZ90nMZmc5/oIlU6ttkWvF4kIgQFNKC
qbMwlyFLGAT9hL48UiwtCC8RNz/Fhzp9gLt3xeV562FLvpVGNBUipORVwQ+S+Dhn
TeIHUb5yOvyboCxpmmVvHaiLUVMhIQzJGrPaM3Wwpe4Yg8lir4Qnr7RPRw5pdmOo
AOWjV+jtUFvmpfF7g36appDPEXrViXb5k7QkI3d3PVAIjiGvB+O4MGmTQEPEgt1L
4zezSvwhPurWVu7cTyGKi/6ni4iaeK+jAuWrAuRjuPWobu8+hEepvGHRo8fccS3B
PnF+hN9uLWsgWTx1ZXYToXm6JazSfwAGd38m1EdzmPMiM3lpIYwnDTTewq0G0nNB
jrbcFEish9VVMBV+UTFp3rB6CZIo6xMuV6jrSH3JE39pICVREuUkjTK2UTbJ1CLf
BLio3oGjoQPSnFjHum7CYrgswqX+UUg+FLCghIZfeNkf3waHorLRGh5rVjOOmKMo
g4E3P2fojvPyZTE1/wy3RebwMyMV+ICsXmA5dnFup8rY31fTOzdTe1XE51wZfmZ8
dL6dPjD6SlMsIAaIJ82EmDIMwIwakgtuHPD+5iyVbPMlqrteHsdAur8rnGthP/Bx
lRdYj1G0PzWUs3y6rOhsh2hnE0GH24cTqiRVx0MxHmirUEBCxAXnTGV1BO60cRZL
oKS/9P9+BV1Ur6H+WDabSHjGBAt+5bbpY+Z+qs3oSMW8wUalXt/4bBJ6prq92Eyl
9tytS0C9jyE3WLT1bxHXPfa3UxJVu9Po6dwwH7r5XJJHGdyk3g/JfttymEyqF/v3
M9zveLGaOQscpkB+TJhGPNWkhSJPY56JesC0Of0RdBKgaOtU9RN8rHc/mwQ2VdPm
N8ACYef/ZHw7+3vIDw1dUrakepel53a2BmELVGvYe1TV43V9HL5ZhFxi34GTAKIx
mSt/O5RWZsJlxqVq+DnJol5V5Pnj1oiUVbvh+4v4qOvTbSt7hcDpmGYfU4YEHDAQ
EnMtdxLGayZeupVE1zCbfPiUbN95s+l3jnMCFz/jbd7TzYsi2zSp9txMprTwNMKy
Ym6vxbpIv5PRJ3kOgy2/SmesfQoY2nRf0xDNUwk3rz0hGfJQX1VtxMbMSGndwSn8
lk2r+8nY2z4hnbvuQbQEiAxi9QZOXiIcCkHI2AJKFQf7ojJXj3utuKiZDcRdM+ul
kFCByOHnV+mgAG6wOFsT2x86W+aHN43zcfdEfHM/oda0m4oB3X+KnZul6T2BcLtn
aY+qdHA5gahbk7k0U1CFi1EPerA/ZtZU7fqGeZCIkpmxwnWJrinzsDb1FBOwDvyy
12DagCjdUO9sxzhrV5hC/7hajY5PMNWzUrNDRTa2zg9Mifep2dwvZztFrQ37O7Mo
Z3d43KFlkeXfc9/HqEKwG4AJWaW2BnCHujbup+AvqclsKDbi3hHX9VBvERcKG+vQ
Qt202oktAFCZx33QF6mZV7/K4P9G9S9AhV30CiibeL50ILeE7E4YZ5ITqluxKWfp
TOfUY41fw+EXDARZ3DPwaC2mo6VqDYeqQrXM/BuElBfkZzLJKa5pDfh/CRo3ga3B
z5QLtcwm3M3ZDFvXqFqUzqwvNxp577s8taFnwgjfJI7WcNmW0DgcS1iull6EZ7yQ
Eb7m68VJOPlf9UlSresYvt6m6Z1DdXqHkRuFNOgjPLLeM2ZrIJi6vXCSrXCPggsm
DclKOVYxsFPwE+Pu3+5XgO9cIX5U4heGd+c5mdIauPCiMQ1QRZVuv4GujidaN6Xj
VmjdVgMPgAkhsuZB/MuKSWmV14oThzwW7MziVnHeJId6hRKZLRIKd8splM8vXbjn
VVIuQZtcFm4dCK4I2FZl8Hm8cHO8Loc0lo8oSq9Wu/8SGrBxhR7IWF4FiSFXX5Mo
TVf5rv9oJBoppEQDT05lgDky9Jfcb6+iNDnpZ7nAH4SpjTxvRAW2s7fyXze2HXVf
5tT+39E2wzSbJ2m9veAQ1QkngY/4OweZj2aDaH85bjmh7LaAxJFrm7DlHwwffn8a
wuHKKfRgf5LpteGXsyLWEeDHBnsIRqK0RU+C3V0qto/06HjcWfABVjXp5IBXURng
Iyjb0NSx8Sb4uGdBP0nQtZOGDG4AX8b0vCPlXaApBuDgx2/252T9MeNfabRGL7ES
0SSDaxrE6ZaTAjswYeX/9q3zs3lhN4zg0pIcsMmmv0LIOfIzt7js52D77i1NbkG0
ILU7/93teKGwFS13SWjxfaURassjomOkymFx1z6t6ASlFbICg2E5RopalhjJDocN
5Oeq50agXZCyNPieZ0F2Q4Gf4EFqRNosL0NlJlIFte/4cjkYAkPNZQebf2yqyPgZ
MCGV8V4ndkGgc1u2gWNRIGVi5BkSzeFEH+RPJYNhYmL7IcTNWir1xQmArq7bfRsO
iWv98e693wlg0tp32WxiAuyQFIOrXhJe+DD2nrDVbJ3mtos5Ukof2iTx4Njm80Y7
PmtYt7gJUaodY8+nd1JMV4/42NbwoVQkpna0DzTYbhOtUR5+pypgyG9ydQQFFxtY
R88s/VudgXTuyfTBV4Rzvoi+YqTjZEYp+mdPeJsdKAB6MlsglGz/0msqpkpTM8Gp
Q8ZPEVcBrejrwk3KojRLL+US2ZUenihH93kVjRC4bI8+4zuNjhqoKf0lChy2rP8Z
/NAvkZHkF0IptSeo89gWfDcbRAtw0ObzMSf1ZcFt/8aGIx7ov+hJBPt8SUDsW9wI
4JaHFyagFq9usCyYXrLki6W4SSM53Oa1/9YI3pM4c0l95DGprkY/LXmxq9478Glt
5+0Bv2njUih5/7zxCnGlvN7xcFI6Wl1x3mmuJAAloKUxWhqbqXkJmGN56cqaqy71
c9zyjjRp99DlQK9vGIKd4X9vb5hwuT06J6Q80SmW7Gu8qLY2NFTFu9RUYxpWgwzr
y2kP32mtAP31+w3XMhV+DNVFaRYw7b0ocpSWFTzDKVcCZmDzTC7NtvPGgI163VZ/
zBggaOOKtjr8PB9PdncEFQ3ZlgYdp9pLT9YLuAZ7+Z9XQJdLZENAg3FSsYvnHDHK
wL4ya1quSxqG30UZXeLydHNXa10LFeYWLfTDnrnDdXluDfTHNBXaZrO1yuf+5U3W
gwdX+4CV6SGX+/odq+2MGE/A3GXWslu0wCFeNhMUhbDuN3w53pc2dc3tTK/QjA2m
PNBb93wpiJsPn64vbuNM1JgPnybmZwac+ed826oMpnco6cU9wVi6TJtk7JolbFUE
2j8No7mhsZJzUM6wC7p8cJWmor8rIphGhaSNjBpm/rwX/Jhkx2PhP1ATL0kqQRyW
rLJLzZreeNQrebYER09IQgbmKphFZOi9zYBx19mhSksyPoFWMoaq1hdvnRAy8cn4
lgVutZN+Wd45WDa5nMoBKUF+pR87g40S/qrkADsT42KiM215x889B3RWpnP82xoA
yK2AJx/U2Q1WAMdHNNdmyIzKP4ToIwrIN0RccwClkZm8wnNKbPzvn8cKUKp+yFJ5
4mfDeGQjN7r1W5s0bFFdAa5RhLW4Z7pMbJf1P76kqxxpWJv0WTEndM9QN1afBhYQ
vR+hONtCY2MVML54U1+RZ/VdBL0j+5RwUnyz/8dZaLxCGdvy1lKT+E8IVDQGGiJ4
dsBmFVq2h7XewydewBuKpeZmueX1pWwbCebng3qoGMnYG2kKCsVwxeirhAqtf36C
rDD6wYexUpqoGclCKF9GWhVN0LJ/X3RNPTGB0HrwosIORSmzHqMr71TCoLKsiqOT
Pcn00c7Nq3KDlNQmbxyt8JYfbWNIQSat5Yi83u8KR4QdH6oPsUdtptu0MmAlekjT
6VBizVmQ9l26pCxteLlnOyihpPC4WUHNuQpE5gZ8FpOvCFbqGDD0f+m/F1ChKYc6
NjOHRQoUwyunS5shTT8M9Xm6L4wA/ACo3RiMm2Ud1dKDMH3qgMq63ZeZMAUU4ISa
D7kxj4iWUK2u1woOJsQW9QoAMrex3Um6Nh9nhhpDQQrg1w4Q743PlzR5qAxtLSOm
4bzIpmZ6UuZspX3m7TnRRF9+EZ4R8CGca4M0jyR3tPVV5frwiV8QKd/+Y3Nw2HuJ
QjNkKsLA1iY3oL+sFJkfGynyw3JXNdTuax8XS96pJfoipk3ZYcr8c7/DXUAih2ET
qYRLNNMFzlsBnTioKwjfhRouZmH27eaQ3J5ky1SrpjAMzmX2Fml87vev6oPrAY0m
ggRbEdN+EGngfrNmpZbH1d36WUnzhvnVgOiL+UFR0AuVxGtitxNZEDRfr38YPKp2
QXXD2YYCj4D/XqgCB9HKRaizpcvqZg1wMXERjkj5OEaC5hg6zxaZnZQfl7zttEFF
xO8psHsdTupXjxYNGpijuaHBu6J2SqT+JZoALnlJsns3Z4tusrl3naofX9KkkWls
wnSWKn0r69iP2q8W8p/xFE6X+pnMHy9I2I4FGhxCQqHiLcGgrRrOXV/joro2rlWd
6ycSI2htfu7gwCvFivKmQDZQ6ZxP1wh3mgK6BVgzrZraYkf+R3LPz8T2e601Xcrc
FWWh/p15mIdvCGkhh4wIgX1OKYGadynuNSIJbbPME6+9iNIGjlO2wb94nxhKEd84
gW21fioSW3kPSiv+kA4gzkmjGq4fCW7JCtjNMpMP6PlOh5Hc1MMZ62vzY3xdM3YJ
CHYsKoZG4eXc2tGiE78FE63KsF3WaSdNRl/4//KTUM7SXDKqa6KaVCE8UCxob5zB
TyDH0ySb3edgAT8/vuUqe/FQitv6AQ7YBG591ILse99C7lBSFjZitwjYE6z6axMF
W7PWZ83qfey3fd87d4SRtKhkV9u3yunyS/G/C5iULEjmhfo21l5yKpt0u8hgjv9a
c7tsP6BXVH4Rg0VW+W4PsOKCDXGYYnY4CZdPzarDg5tXdA0VEs6RRpl9n2n5SiwC
TODRbHcW0KRQ6FCl9sLw/4G2EbtenZ8PjnhRNyzP+eta1g4WCJR567o3FNwoRpri
PeHpzp0vn9pKUB1FrLxxEMUkMAORWHbwFiw2e14EHj5Z4k3x4VsnYDj5GCBYSmoS
R2mOJ+jTg+mC7/o0MPm/yrYdwBoTc1rpX2w9+UlMwkuwkcAs6CyrYepNfhXb1aDW
dBuMEASnzym9mXMPvHP1a84qst1QKjzmtCmRf6dMmuiW20Nueyy/JUjSSRKDaSuo
UBDQjxP2VXGjS06mgEDhcsnjz/Z+4Vpc5/bQwxnQXIA6DPJIR9AlCoWGjjGprNKu
Q3FGzHia3CFB/9zvXutkXTve5Pz7bc0lQtgS7TFz/hdfcNVaGA2yImWcgmJGCjKv
ZoJkIM1dXSXGSvp2eEEhUnopiAsuTfyLQA+FhNezreijt/HJ+sN2Hay9F4G1gCpc
eeusxtptFy/ksEK9os8ToGJUQ6rLf/l2iKEd7hjVgYOOkrRwcmt8Vcm40i0BEDhr
W7Jchis8I4I5TwDYFGrgIyY0ZY+34/N270IVUjjUlbNw2ViB7KQ/nDJrGimaL67V
uRxFklRCjZIFkYLkKUbhw+HLgOEsQkp1o5UuRH5qQJwj0oSrCe+zl6UcUDYWK8BC
tS5czoXoYhBAQYplk0qzeDXjvEe910eJkV3Tg2xN65yt2HrQp68Y8KSxQz1Ds19l
xgpW3ciH7scnivoQEMuHMZMXz+shi2ut2y/alYg+rWgFyVwPFr4o1E3uWV5pBKVa
+FF2HQCXq0hMgNCGKb1/zADEokrmyBB1IRrpgFscCsJ2nnllcmkFrV59Y1XTcd29
sHjvjx0C6JqWujTq7xBhCoex6tsmQConvuVa0gzkLRFKch1UKyMRenZelo5hm2AF
Te6E2oH9IWDp+O6CDn42vZcEUo6wCrj4qcx25OHUeDp7SoEen+B6pTIbWnXsGxVu
h44vneJX1qKvkmAOPmDEVkHBB7yYm0eMhGok+qsHptJKQA/GNfhsb1lSXZm0wX47
FF4IGZbf5Z/MXpLoxeVA4UGi0YQ62/ahdfU9Th/99AL56O5WFLDceLWjLRpJlcaQ
lfLYtvy2Hf+zLbiEFL+3PxjEVb+z401166xwBzERvh+iUOSH2wLDCIpJz3UozdJ0
mAlXyPKn/jAkJpRx9MgvrsqEXAajcFCYfJbM9aRrJqi0h/tM2/q3AoPs94JOx9Pp
cI4f1jIK1dZDLEfE5JVISLeS/XtlqgOZDz4gRWPJwHq+aw5bkCI+HArYwd60g/Q4
wOAYuh4zIGMwKXgdOJJRZkEYxXNznqu5nQmPJnY1jWxpL1SpjtzQ33coJUXQCI+0
AUoS8JnpQnfoBguQrMR+RRucppBWyV9//XgEzDUqZlfUF8xqP2e3ZQxNkTigD22x
WzDp3GLNVujj3gSZRGpjyi1lzW0029JOAgvM05Osl3cfM1kt+6c27hL4ElTb5Uyx
vHvWTxM//Lvzm9eYUTeOJ7dwoc8AqJzv084Qb0dJH4kJZw8+T3n/bJEaSJ9uSYne
uKVeGSIkZlyCMzPT8vk3uKJKBEoZtMfi5d3C+Yh6XzF6fdlgcjztvPzEvmnab3uN
0vnHaZs+FA8o0+cmfCOmD4G2yPmy22K6COY8SpFxOneCOlQt/e1FAi1WptIeExmx
urzTbvE4zkwsdWPCu6jARcoRevhysASfiZ7sWOY2Wz/wmFz9DBjRIKu62L4sZNaw
GZqzEx8rEYxcZWyEi3w4LuNN1EAA83YpeIxYc0OGN6QDPVqj8panOpBvhvw8HW9I
01b23bGPIHe41C7w1RGzyppm7P3EzIMMXoiS3iciurDGAR2+jPsye2WPlvvjLx5F
7w76rA5vs8adc9GBma0bw/9feBziO+K8jA6NiKIORSWQSJgKBo8Pzuw7LwlpYSpy
/3kVkP9hZrRDJ0DEmqIaQgwrxJ2Lw36WP2ajDTn8UdJjD1C5ry1eHe/FTB3T49RD
v6jCQ8WxEv21fzEUA57ahtpQYB2KvS3wStVIzTgrdjJ92Wc3y3pM7a4StNHhsEA2
2Rr8zFSLcOtZOz7wz+V2/uM69IKc7DCOTM+YZNRR9hzmnoYH3+Op1axuoHZ/KTJf
RA1BVIY3z4VYXr1M9mb9v9J+ydqYXORS36iiH4eODmmZ8U7JMAM9txTpKPrkm8xj
HsOFET0YAB8VzIpzxMp8vv2fbJGwMf9tJhOhzCH5LVfftXrGN9OlnyA7E8+wRcwA
9bdi5cTUpqmUc9D9mxpnqP8nsRp6e1QSoFcJ2Of4fTwmAs9Tg3qz8Y+0/9CA/b5h
MPea6pop9eGQuqezN6WqzhQw24u6Hr4y59eGxzftmv7Qdt623PpbJapKltvhTgXa
n73fnexMAr1hp0j1RDq8nWyty2+SSxNgUHrbpJl7U0QizQPBiFZa7SXOLEES4TmZ
Ogdlemg/l428+eOitFU8eg3DAqtjhRUvkMj/B8oecoVlAIlZJvreOW077WjU7VSr
xA0PWvEfaijb7r7tAAlicwrkN6aqr6PyHQ7AJi/Nnai56Ys0/BA04fH9J07F/Ut6
SnGHbwr8FIvyeX3RHZZCzOVXVI+/q7PuoOiy4mxd8EX6G/skEb2nVp/0Jwy0GUqE
eV9kw6IJ5JbCLVik1rAV43vvEJA5C+7JLDRCQy8mkItmsa2usKnwxgssyxDKk64d
IAwxToEumCxsPd3TB+v8+r8pCgiOGMZcjPN1x5fM7lgxB7Xx3psBqg0I0fcpI/8j
GtZGr8iSgov6gjWi0iUp5xX/rYkmgzcIZn6gmcMlRM7FXcrFMCjGZOVnQqfjMZXN
hQAeIzLpP3nIa+5h3o7Ey1s02RhXDu2Vg4zzmYsgNhrhuAkRcEDKWkAi1+nioxtR
GbxEIzkYUEqBqg047rY6WZ9EtjTAY/EhEuaVuPp4Pem63Hn+BP7+TNPVnlhbR78F
vVSj/EanMlpaHReXNmZterBjqQxlYteGqjhkYhWpPdzHort+8dRz39yX4lyfIg5+
BvHYA5M1LviJEmQP4caXf5pZk/bJhJjyv9pHj5AdrKD1sNtrAIc9cPIKd3RxWnK7
9ER5LDeToEQI4hHY/JqxugBodjRqNJeQ/Ca4SKWJp5Bu74H7LhMhsHmTY+RbqeN8
aFWTCAz6d5Y/od5P5F9wzIU9Qr5MD2cHN3EQrxiMALee073PXaILF3UcW7DaR8ri
q3baSbgv7O4s48KWRY4BrTXxpx9Rrpuh1YpYqX8ia9Us/+EoOuK7N8A4cm9glOky
y5Rr0GO90XS3Cgnt18wIY6c/71NGoKWM3R1SpaO4fMYJAep/Cw5tH65ouNvQoIg/
GSLgJqKCbAlS3E6BQ6QlL1pnOr8tyNxtLNIC/q3g5+r7IOkfev+oshEa2BnLsC0B
42G05udIvXXFmmYGBjFm1kCtrwe2dXKneZ0dfUL5Y9uWg1V7SkNK/EzffVL+OM0A
A/yd6+GFJzBngfgykYh/vVG6A6aD7MncnpZ8//g5mHtfHRRpaDLxFcUUje3H+Kgu
hWMXfHlSDFqGLHj9v01eH9kOCmoeczksAuctMqh0BReR9bGunz91KvW8Of4oynlx
HYp6EMSPFLdmceGougcyLNS/HGfrLB1jZmvgb/IOYQB47YPTIqlJbfx2ph3tvGdl
EgtbI9L0RSx/uoN9dFiUgf0peVCt4q6reFPmokDkZ3gbGc1rr2WF0ajO8McQ1oA8
qM9uQAtaOQyXhtJJWBdCGPZ1iT7sHnFoBrLHBucxybiZ0GZsuVXta3ENCbWvLCS8
wrdKVzWgQ114WUO/X3/dqW2wUxY1UU+0FzAVzr897IDKF/b9JxzQ4JF/DhFt4pF+
nIE1Xq/Ou3evKn+/hNz7E4NuRHhm+szJNcSbFthXLGxgiI+eoi6llaA7leBfdVFM
75/wksLgfT6rrmIo23n4scAZrWU7N/b1wU/nwzIpltXheAWgCq4gCqrsQ9vDkupi
jRmlapb1DQVDU9koKgImVFAndj++OEOBDrnYGtv1rnXAF3RSFISNp76HU1BU1job
bvlA+nAg65yvMOiiritOXQvdI1rrnqDK36ddrz9pcUcpoFEOWKbcUrgK5oDOUnyq
eTRjajhovPn9DQY3YkIdioMQ4xp54yAgfJdKrdGimPpXBKX+wzdfQIGV6OKmXv+E
HMdhcr6GK4ie8Jf8v1R1ujjFSd+pNRUEUNTMPH3ma0jSxOnIH9CmSbWaGirYNExV
V60m6hD5gyM11JGESw2KxnZPptfDaPJSR79HEElWmdA4JHF7AgeU5+fxpHQteOX+
wF45nlCbX95Nkc4nmp5OxyB8BKLrvBUIqhUjHzsFhTFgpJO+NhjgSYtbxnWZp+uc
FxiXhxgAPv0jOr0BdO5kLmWxtAe0eqjyHJqFLnyk8PYmCcPGJZ4wfTTaMuVicTzj
4ePYY0KXdPfjnntPmwfx2+mThaAgctZIRhjZiyQvrxPPlzlknGbZW+WpOIN9BKr9
C4EYjI+QB19fyhCqC4kN5pvDnxD881KzSe7OGMB86dipJmBweKzDtP+YcjclDyYu
j6oD5naDg//smFb7r5EwXlOTEjJzmT3etHkrlwYYL32y9b9KSJTMy5PAIxcl5LtK
NrQ0qEh4LASR9Qg0xa5FMtDJpvJw4TYafr8c3eMS/l05JdbxZ/IAGiN9NINhmIQ3
B46i1tlsUWpCYmgotxTBNkZJ2uMHCQx1Yms+VH9ScUvkEZ19h6JssL86d77zhy4/
0McPHFG/g0o7+bLWmM4rKfWaTyfBSfS4QUZPvB8lYb2yX1v5tzD4Pa0ovZJbFTFF
HGwXbwSx2mdho8+2WFCT5PP2sjQB5uJLVHsiljdxE9TUR6dVa5/zmFAicRzr6XMk
If+8BJuB43UeRLS0TYQwtDrsHHzbvB6LKKFYtYexoXXFVIn+0NIf3LO532PvapMk
XsZdA7PnF1CkBbrMJtTjpS3XoDPsRGWntrEZWVIe+6n7UCaMUsixcL0HQoCFqTOw
hcFREWSjipOkeEFpb5F22vcY+CwQ4uoMEP3IjVBWzxQT3aRaDC1OkDZhMdu42wB3
88fzpR0gliMTFXV/gCRS7Ha1B3zolWPHyuZ+2dMFAlQO5qNTZxniJJAObXKWngYe
DuigeeMomChn25XD5VyvlQF7o+eRaaH+qOmLNrOlT38HfUwvd2FiklQsqq9ue6aq
eSAsZJJauTnnNT6HgF58jUJVXlyxYrO4umZrXD1uRqjf4boAcIWeG3Vk9jhqCuPN
0PeudGpOZJaf9uM6UBwUW5KSILjIGBtr4jUAQTp5d4TkLVmezuP6i/UkulkZ0Jhz
900KbrgEfLq6b01HpA+G6XvOhe4ButTxiBOWhIQl6h8+hCbCwSGrXW0ZLsWI9lRE
OVPcXjmnadCA0t3S9AQxiMFEVn8l0UOv/Q9GHV2KIw3JltTpEXTMznDH2yhbvbLk
3hmhXzJLgBn1nA6BNgQmroUSLnptd4xBybqpOGCvgXY5ajzMVtc1jdpkH0plsHkH
MDOAe6li5vrZ7FdK1VFUX4QceD6k5aZlEJkLWHip0LDnoonYrFHK1o0dEpFeBzGn
98FIFHJo30Y6IzroCWOEUaJbpCqit3Cd9yejE3hB3KdXPu0cHDFwXsOAunIPlBMq
TJBI6KeeDnJs1U+sR4x/lmhBx4p6cgvjaqPMqzWZRMqQVNERx4hL50Vgjk333c1F
y/s23YfqER8f8VPjMkHzoHE2SV5Vl5QS51tXyChMWTqEs5xzTvhnxnWfwusVJbP5
9dS5E6FsOsFsDGm0uh4rcq+/qFFBfeBfShUDHk0REQjXU1ptNM5/ShB9kEBkpM9Q
j1NdIZIiAMgRquRYFpHuRWgemU0qZS3xVv4sXN1nJx0GzkQgPZvf6P6EeSxfefA6
zjAh++582t+/4m7inAk+NrCrQvohjsjS/Yyom/koh8nsjuvHpxz7wCY8eCfGQtd4
IGWz0no4UeBx2lWwzeM1xdmSfutzHhM0UMymQhelgtTXgE7KKIw1eGY1pCPXVkML
oalCJi9sbnPM6c072DVfsiyn40NuWavQGzlJLrfIJOpxjDAVMwpEv3WjvMxb/TxR
sjxsaD8BEjVxpBz8K+kCTuVBomjxipUl8wrdwBbKKdGYEFpipmQs1a5LUGCbjj1m
oNnTcAT2hfTCDeD9petnmBt/iGdClDgKHLR7OtozykQBDJPOxXsGyNngvqU5cpbS
d7xIXNtluuAEs4MMYS6hOSjd8ZoAYpR8GM6CGHzxMwZ/Wq02dR9SW/kQ5Ix0eX8c
h7eiB0du7t4NFYrmj4dRhuT8p2Vl9TwI4K4PeMxgaW5ydVTopUWlwoNohfutnT4J
kuoaf6Pi12YkTFICjPK9TMBDkbCGBorajR8P6E1ym142RytnT6ag4aV6QSEZnT9O
VIYaMTP66dpsPHiIthDsjdwQGnHaKc7C3vEk2dn9hVQF8P3D0npwmzk6DMajLmzx
N7bhqFm2+LUYneZMOm1xouK2abR6ttQ2KJxuCmyHyXDPWOMp5UBjh6KKBNmFnjY7
a5xAyQ6CUWk1SHu5ROVLtUvTvbeHOC4B7Pj9QP8PEMbn8V2cLmF+PD5BCtZPfUgY
uyqo6pu1pIB2VWZD6bI2e7Ww6219/Ti5cAVmmQVKCEmwsKPO8x0a1MJcDc53lRRq
dRI8z53KKLbmpXXzuwUFhJ6IEGR/eB4C5vrz7F/1aDgWwNAJvH+JLBv6YCtdw1oz
0jabtGFBtMptb7QGfI68O4rvqT9Rz8Lvqns9c1dVGmHvPLIpx7ZK+of18V1btxPd
zShak7NOtXpqvNt1LQhol8y4eX04DkyHF1tiMY+Zzwn3xUSRUWhG++cIJHk79NqE
vOOotQKJtclBuX4shf71WX6L+9CnCcalRDd8XKJ8wKCGMVwzT8wmCC4taubbdeuG
s8pRiEGD3zJNU13jJawcF7AaOnMWW4G6EUkGGc+LJc5XbDssinrNlFCAxprSPhU+
VOysiGVD0kvr/hfYcmyrpJQnyVnGE1MC3ES5N7ZCOpJXwHd4mu8erGQjFYLGywcs
x2/rzrI61CslTw/ohVT5QvJ0HRhEoWb0dHfhTQc/2N2cCEqFKJsIW1oINgN35h/5
Kw8Bqmu0Xkg8PFeLOzxYJMwXl278UR3lw37xR1L341eMmQnVQfakY/T4G2eNqY4s
4Oc/mtEeJiWb8UvZ8JRwV9f9nqSowZdBlnjq1jItT57FRNsU4YJbAbT9ypTIUl7D
1KwQgNgB0JYiFJnBRPKA4lVcOF3Em6KLiDn0XYPdDWlV4/vHd+UDu2TFagybzKYp
CCaVwkUoId3EU4Ur8qFPtsFM8DVfqbmK7SelgVYVE+46s/dWWWMc5UxMQxVzFTfV
fTWhjuOYhk1xc8oRvQO1Ij5nnvT2F0UxByDaHZimdNg9uH/L8CBPbw7WXWH19GsD
ztJbPSMFDp/fzN065OMSlVyyTnJQkie3AaKrmnHGiF1WgOaX23jyhOb08sN5O/NZ
mapldVJgODNGVMOKEoK+zURVV1AYSCUoIr2YZ3yPkME2AWcyu1yvDrmWckkbOxLW
By8XiWRTIh8KHPasxpsBBoaHmc/pi/1+4RZ8FmPocjlpcAinBQMa6qaQmQ+nygL/
GRktd0Hkh4eSWNXpk6uL2HFZK4eohqUEvM6T1BAgLqwj9LfkpEnlgv6P03zOyIL1
7DIm6ptfFpj6mjdEyIYvJGgSiUJqs7/NrAAWBcXI8opWM4i4aU5+RR/hM+l0yYL5
By7q+9Qjs4DnAXwWqaeWJnf2nkWw4yXpZiggRluFkjuobHlnK/pCcOL4TMOQBg+F
zufDMnqbmp1UjyTm+Jfsf0lqsTTNtQQQRaLB3uOtIypG8nI4YeXBLdsAsy3VsDnJ
0jkR0yGs+5h49kyjMn6ValrxaRQCmSR5YJHDIZnELhJODP049y9FhpBhf+KOl78n
vEj9oB9sqcis/etlnZEKUpnAq8WcP0ZuGqS0TkPiK6TNs1zpWBNjrTgY5Tf+ZQO/
SDtzwa1UNJQhcKM5Ch4llzQUGeEjY9yJwU259sZTmh3fpO1Zm8JU2IX0OHZ+N2Yx
epe4ZDpAkH/30IeW/wif/aHm8xSkI2IHX4m0IbCjFeMp3b2BlCpAeInO/BTKxCSi
yez2+jDIZUHU1NX6g/4iIO4aMBirZCT9ie3UU+zEg1CHd4tSOcYCDbOGGsfxaOB0
Igl9RXAW9u59L4KB7lX06TY2+fHWfXiV1h9eUoytvAkcvTJ139lXTWQ2yTqA5A01
GPC4oaC8xEdswnWKcFWvYmZ0CalHueNz2nxlsaRl0tpXoLmiA7IHuhx3WbQwZ+Af
v0xzf4hjp0P52oMjqubhEVV/mIFPZd5DRryt6/OAmsj/fACz4wKvHYoHSx9Hkkmy
rkYWBBwg4ryMmLgk83ynjuf7arQLGzVVwzB7LSv5Y6mJBcpGX4fZcbjZLk1KdWr6
MNyTB5RHcECsp30Sz7FOvrxFHWB7W1Vj55QOmoOPEQlcG+5oH6iR9dxrexiGpo92
c0Zrcpb2NG0oCuMtqm2Zf+KCJMgMZQIvboqChkruWNRW2jPWGiR7AguPXbA769uZ
aCGHN7+TAtrQXuPUdsC8+6NbgMlioyUcKPjpCio3go5Qy/WJWCVKbDmgja8imFTM
ynygC6VpzcrU7a8404NlWpzF+JURI0OcQTQifm89ghjYQszYtD9lS42iidWeGnm/
Ic2S19F5Vf/+cqESvg9tWWAz3uokpbiObL+EieXwLjlsHWBUQYV4WutHMO1aQGLQ
mW0Z0lUAEzkDz+u6II9jJXBr77vAHnokhLEhNne7vhS+1wrl4j3Poh4z1bwehJgn
EKINWjkj0SVriSPVJyAJ/xhiAluyv251cgYHAjW6jWi2Szhq7HZ+VJ0pGU8JScsd
SPadkszt/OCxAsR8zC3C5wzwfTZxiPeRDPW6oPXqOSkiqRf25bTlakaQuTuJGnB9
m9cc08sL3JhTnp/4wqcgvor3BTmGcGHm7qTM4wHuYF6wLuXuTXRR2UHuNx8sw7On
cnlxsNp071eYpdQ7yZJm7llT2wH6AvXF3+2XljQMFvua86606hboVcw4EJjdvy5+
zJbwmohiDev1RPYnj8khfXgB1fnXvMjSEN/3t5T9UP5C+O1znrF9CXUrTavoHBvO
TA35p+G+Ie0l+g05MPfQamin+CIa03WrIsS0uEGYpzAmgMha0NK9DuqZvfgu3BBq
we6jdkBFrhKETyiarbpb89fAjKzCJr9IvDVmZakcdt0zkNzxaNDnq2xmz1J4q8UR
vWDwQUIA+oZ/D16O7CXYFYGuZcGYoZkC5IhZedZpdafEAnXMXQo+QdQ6Lxx4Aadb
9ciHPKhRMCK38r4y0TAsErSpxX0trnu5gBhF0rvsK2272yAcDWPZscLz4yBk8Jai
0jfrr6qo/Acg2z5dhaQfXSQYFwZ2puGqrotUpQ4+aqP+dufL2BVXFR/wQ4hOH3EI
iyC2y8fJS/U9F6AvVFWSNuGzviuDvvlM5BQbe9mOU7uuSlR8M1qaK3c1RRR/bEGh
GrHEdS2+n+3pQrJbNsER1SbvwglHEpiU1icGqB/9WfBjBpv6INk0XZV0ak+OzO1V
w7qbtWY+qTJF8kyG7LdP+WJcQUnOTgPLqQg/4fPOC1Pqu4RQ5suC/QSP2r8fJgsF
J2NkmiWZrik2hG6fRDHYaLc2hq5O8IwDM2jIe7LqJYp/CQ/C7b8R7Ti4oMq8zQFK
nvkAkToKWWPt0qmVwI250cPtDeftjDz8VG1qdupCIol/Xfxcw8Xt3idlIc9kBk4D
rRdzGm19cPWtd0jsbdPkpqMRh0fpzaXW5d4BgkR/Xm4tQEm86FT3PlJk5ry9hAFc
EuuGXF43/KbDXN8aoDwLc9Wi2ebOjjzbNhT8yR6E6MDgXg9BXn9l1X2drac/kvSl
fnf69pDl5jlnFCKmx/yu6Boo0gmgvQ2dmYp4cEIhYr4NvFh1qZ7jStmpEp+K97V6
XD94abiWq2+GAMNBZPtKfxuIw3JwAJLO545AR71gRZTABAqLwjmuDQgy38AjoD+m
N+tbOPrndfl3Va+EqqhndjeEmQpHMjtxOukCcbhgbfPzpqxmPvMBb5MyTdx7RUYh
yy0i1f4Q850S/geNHdtP1/qqYN64w+1BBjF8O9QvpXUQH1i4rgQ/siv8xY1YWm9a
ococQvp0NHCnFrfBSQhnkMmCt3FBR7r3c+0Ct3AvjHWCECBMZaWlVLOoFZ5CM4Sr
E2aG8DD36RbaFu9DRNLb8f990VkM1rYHklSNv2yumL9YjhizkeR9KuAh+YJvFmoS
OjU60iW3L4igsxUGPeaZ2uRZiSOMml3v+IvA2Os5YBoPYBiDq/FovTpRSMw0LMPO
/y2Ptp0jHWpe50vSTQ1AX0c3osOalmbbTEJWRG9DM8uI2LDkaiL2XYDMF0ObkosI
vIkmr3VtzgUgaET6lb3Trn6Lc67Bx/Op0cONc+h5GcSO05t3kpIDj41ziZ+L86Xs
sQ0nwaZ77uIM5wFVum9ffeKWIiaPpyIet7u0aY35EM4I/f4UbjSU+1AufY/b7dhQ
rYVDWyK9owDASLIcX2+Qs7BM2MvpPOcyzVARrPRqMlFmcKrs92thcNs2do1+t85j
bLB15FOJ66PikitZb1q1Yb02R/OkjG0hocEakqqXT8WIjAqDx1vbdE+gdFk8IEmM
daFz7XBx2xu+NcZ5Xwhizab96Tncq23nKhJe8Gj52Qeg7s3KFhv1FKlI+N0P4tpI
yS7y7nKSr9KrGGNX9M6xRbqZw02Hw/iVttjZ38gHBlLwWYwZ1dUQGQxCQ9ytAAx4
S6/fy7BLvtwbj/W7M2qPR1aVDDOFYU6+hfO7sv8zLudCUdqg6kHVahQznNURk/LI
61Kvdwu5sFhfGyiXMUozxNK4qFWlvLOWx/jIxduEPWaYgzemg8sry7s4bTacvEq2
7rBv1ymRAJiP39joVkqwJdmEPXy3ok+zHEoSur8Sy11tpQ5zqma92wC/bR4cFTgb
znaSxgfvmfJDxBQumvjQpSTn7n7APd9YZ3Sx/mxSPXHofU11/zLlnDKSd7xqTwJ7
Hlc4MAOpMVwHmj+mOndph9ybF/vCs9AbaB6gZsCmQTe7moQMB1sfJC4MZV62JZmT
sk8z/ldlJzEOlmEsPC5eRa74bYRx6vAJ2lfS5IrZNmySHjaZUJ56g4qDzOBfz6fn
pbK+1zWFQhBxvYsHZBJKIYnkbywXAKESuvIuw3l6dO2y+O76iR3b1dF9bm1KVpyw
OpktuyBUHQ1Wl2RzQWqOYlNA5zo5/ph5C8bwulUU7APzMVADQ5wgwCliYDiOxRYu
M6AYrj88OAnwUjoRImtls/rwM4KAAvh+T0ZmqDEJCRDRR58crphvBAmMwD7YElJz
h00B4ykREnJlKwl/1sAm0ox6IUQzWZqKHIRV+7gOEyYtIoZxvVINS9TKHUXcPqhV
rd0YgxR5tAvVTAYGQucusjRfU9ZS2rqsp1g26Fbf2zI8wg0RVuE863x22gqIEHvg
qqqhDARl3iGcSoO+nTC0AlhP8BkppFxWYt6p/7e+tS9qwxHFWDfs+cf71+a1+tbC
9zMH1rf56CnbLGHes8DeQnHShGkFTVzNT1aL8PqbOQUhS/WK+eRNrcRBFkePiT1v
BjEIZG8Z4NrfZhVikhE3PPeFTkJQYkjAfoFaDJMjC9/fBB423vFkXwvg8DzvWTvn
KEVGR0oUDW3mzs+dkt9qoD4+LJKO+GIxQv5S/LQ9DY2/UDrvbQpPzT2ovgrQMG3R
iZAqUNycLWC4JevHBS/yJw8YCYFnACn7xcsFNCrKnreD9l7IJYLVBeym7yu7MG5I
0LmdEw9CTiWCWDSFZMSrGZtsT7XlxFcaRAypHArwT3hL+A39OVm6Lia0KSeqJPTu
oz9g+m73ZTTxC0oJlkhNLuA24bUFra5GodTqzn/3Hep99onZKrOHo/+TI54twLvV
EiOVTVU/U0I3MI3pkkHMnfGOCA1XZ1y1vrArLknH6JkBY7AWGULmK/g4Wzwmz5oU
XNczzsrC4FIN5NFHjw7TpUPpfLV/MwNKIoCXTAxiiNJQw7YaaAai5whM5tnfmq3n
KbC4HETW85LJRAuBSNMbFrtTPL1HWfZXu56/Vn0/sMG7dh3cZATNCeDWpIFUT1ys
ceTu3zkUP/VPRf74CpgT3h/aFlLMfTjhmS+vN4wtEbG9HrUsGtYSEIE5lSFBpP8u
QUCsuA/cQ66aBnN+4iuX6F+cxD4/zAc0omD9aOhbgfVWIfqs8c0KRgcEyHYmIE8D
UMXptwu+i8T2BY9aSzKCRDQfe2lIXHj45Xq/0o7HBMbnCsLVUZfy6T6gAunpnDup
hV8QjAuIgvKJWNrYhvYmHd8f6dCH6jm1FEqsl5wjH2rfxUwE8e+Ftr0P5wRSB8i+
aaYtLI3G5xdDHxE7pvyK3o18f8i1qC3wDGcJ8v9fBOPlUi9u7iRrQgflbl7VLOmx
lEbPEt2KwqBOj7o2+cgB/dfkRRQgJRoFQAdXO0mJuthH81wh8loHWz5qx0t7jr/T
a1Q2e3lV5gvUp2cUWsyp/zVmE+oi9BEEaIygkQgFi6pgDl/bkNene8HOp2YTE3Gm
bTEKbp6ZHNJ29xLMm0LpBVOEBv16KPzvpFhVZi5OWIrKdc0k00dZQ2zoTM5MSJNB
rqIbLC4A7uXeI6hIudeGN0yQoP/pORtR4yrCjPdYRANKgvawg3EH1E4PM7rYj834
/1y/qi7a1AESdydcfI4Pnd7zOgehIFZ/y93a3afM7upMFgPvpl6a5ew3KRYcqgx+
HITerb2rmo/DHHJD0bcTdT6nduY7mhgsg06T0Fs3MCimA6CVnbBHu8gIrcQCzBuS
t35XOCVZddeuPyeSFE0bAN9FMiRfbfH3cQF1sP2NSHlSMFrhbwQH/zuEcGqtUWCM
WlL0tEsugiWjRzcTKcgieOvpi5oYFVVZ8/YDCYo/obOLPS5JQAwIBCpOq1FEw2Qb
1MZGHthCfjOHjuimX7sefmXOQUp7kf5jSU5GLKdBA7+7kbrYZSrHC9z3Ay9tq3Ce
AUGmRhd0SsbIlVV0lbFGxSeKmgTfrEqNibKJyh+FSjvFMu9S+CF4wZJcYSVwivJV
peqpqwWcpPDJKuxOy7bHhkq3rV8nmcqcDjck3MxJUcV9oMa008aUU1VgtWXttlaw
ASSUWm8jachJhhE7KLQi7SeMbcpFN6tgy+gNMyERm6ut3JiiHH2UFeQ3LLiB9KzE
GCTrZGwb9JGyS2iDBt+fPZJUmya5DLP+woVJCSHQBrjm60zOkrLV48EUX9oXfoBD
uJI0rijFq8+pAJWyX21/+6iQJjXUVc6UcitgZLl5Y0xdYlmLBwWL85V4kJtaJZub
eipJJ7XYlNzWzoTaTLsbbFgKEffM3X1toj5vT/6fRcWv8ejT1EhnMzxGBNmZBeQk
vs/eT2wHYUeILybGMU2S9eKG96hIFvzUn8j3HQ8aiQ7ctKsCl/KuCH/yiSZN7/tn
D55hezxbuMxNTWp0evfaDmZj1Z+LpDj1IGCHkOfmlX6hIJSmSg2tb4gkuS8vHTmK
P+J3I0mFkr7ILK5bbBMFKXlmJS1HpVim4SOEk/430KiuXGhwviVWzjiG1VAGHMQr
4DAo85TD+P5xZEaix6c0tD10iMpH/kKhYMqK7nAZis5YR4/hawgWo2EDT0FAeghz
AWJ5F+jI3Go+tWt4qxaHfiH34WvRKFjjtrxSRTXTqft3Sbgds6wGLNpCZXK0ReXB
pTJypXNyDD/JxhjO20beJmGxKH5OMe3AcHtvQCSzyni4McqLzaRSpB0rLD+8N45/
tVmK8yOyUxRG/oFUe3LlPiQpJRNUQ8bRKfvyTtnBtVGT4XB50sTsfiESLHHj/1Hc
P3G2RxPPIewsgiu3byZIywa/JBP5TvhW7ViCcZd7asYh08BV8jJ3K7d15W0spK4N
9NIGQ9IjSBgmKurCDLos1xYoQCrUZdRAdBzbuFggWwW+7XYFiJsqDLiBTShmmm/D
IvH1RM2lXqk0zHi2ae9ieGXGWhWXZqpzc1al6uGbKJww4RrwsAXzmkhs2J1cF/kU
84TfyfB2LLQ71d/f10BNg2/FmeIBM0z/eFVY1gG4c2/VoIggupRRNaKTwW1MF964
dSUEjbFAhZBRvE9WbISqf2X+uTB791qkQHK1mGjxEs+SI0NWPT4s3Azmn3OAWbmX
804CwiaAciF5B7rj+6ynWNmFxGqFFnrtSkT/6jF6tVfufbjt6MzcyDlL5bBe4n3z
UVWEqABsAWytRKuYRVua4vsdyShKCAv8HgP+5AnXspcveUOERAXbkug3ZrAPb99I
MImPmp6Vy3xe141SNcA1bZHKPpCMGPPZz+yi0qrkkRIQ1T5W+q0mwjXN/r1Ee7+A
zwtTY9ZYwlZa99R75ciiwK94O9Mbdue4IaBzUPYTdUI3l7WQzPIL5OOta11Oi/8L
bmAymwtN57LRS6yBJ3H9i6300/XJWeYpdYXm+w0njiEA9Qxv+TGwzfb6vUh/6tNe
jRD3ZQqRvgLnfOtTuspe4cNhtoGFCsAZIxZ67/XMjEy+NtCSvxrxlX7ugfON03Sj
ha8mhepENM9JiwduVnNKCFSdByykhlE85Nab8JiThCFUSjJvZ8XBSzroomz0kMnr
rhyIz0Uhx3P5fLORqrD1rfe6VrkIddUU76yKnAgu76A/5ZnxIhuCIfrayMznZ0nV
67ZtDlZY5dNXlR68HMm3dU+iVGsS+yJ9bFnsj3SwGFK7YtuLtNJAtZTfB5LecKJf
rd5kNGi/ftJ/Ry8SNtJ/83T1P6QdQTc/2eEib+n6Lm0iQEymnqf5mWEifAlWctKp
QcKqgape1qecmw1jmI6Y/q95sqbG0ink4Lrd5YZDrtUdGEJaMUqW608GY2YhFO4W
cIZq48cxPNNlax2kDTAp9Ty/OifpoBcUEQglXscGDq2fos+rMLcsfSCcGqcOFUBx
odC4gaCZlMwLSrxrtC+4a+cRiqwn/uX2H369MnhCQwy9zqTxd7qeTZbFuKnf7aUO
GSRHKYtMib49yMwzacZ1RrPdBAgFMDWVhC45C1R5LBgdMPnqdshwGGc0puDDBsj5
OhD3sZZYZLZjFiAPj2a/RtgIcHLL79zmBKWlt75n6mTOqsoGaMxp7QogLntQX7TQ
8A3KDdZdEK2PZ0SZP9WYwOcnKRU2654EWGjHm8+vLKhbotJ1SFSCDktNkrtKMkgJ
94FHguV1XWg9FcTngjulappzrHUFdf5Ehu59dIyT5k7p4DV5XfwP+COLXsXzeOPP
eqtIJWqovCStinlXpWe6X3X1p5mXnMUP8aGIBVerABlB6I4hh6JBTSUseS02MbIL
CSI/tB1WEZb7pcmG0XEgtVouaU1J4qigEmQnAFCR/S8Xx35GtDnmbiX/iynwZhvf
6wuT/aXUUc6PUFujQncYIbJZCo5iQFVqZ/PHXZ6sEU0SGNUQ1D2JAxXxRZETXEtH
5yg2NwQOZPJrwhUFA6txNQhlQ/2fi9Mn/BjRli2L4BBGHew5Y/o+zHRsK26zCwt+
duq/NkTK1c3SrtAIjx16tVWWIwCmF4MGShimIkfzKp6d9T9EGmS1pUonozDUngBW
vLPNiJkCNakZjFBLnCMpDOU8ePXRjUuN/zDceb/LiOXwQM/uUo4B71B0hEv+zTOL
ZIvX7Iuc8Qx0hUyc7L/8oOEbV0Mx1n62wf+6U8emdN+V1cB6PExk6yGlDMHa7iYL
Fubdg8Rp1kVT5oZx1RPNciKanDS8JxUT9MXgs+DgOuVhkZU6Ff2Z7kcB0oL560mP
WBhrMgj2B5HGYlPlSY0YjZ7PPEcPBSQ8g83vbJl8KQ+0+GJbUvuRC3ABLogECZSn
yNuZENebAyRWSYA9l+6trpwef7AnpTaZMY9apFzHcd0BZ1UZ3glWJlKtkfn1tU4h
XDM6wv/gnHnrr9sCqdr/ODAAe5Uz9CwomqURBgUgwLCSmkdktRy2LjRpW1MHE+7L
IATNIzx9xnuCQzzSOV9GOubbBwUKY59wmgHbFuuhPXqjvMF2MunMx4rUniCSyo+U
8ya5UUPW+apdXWocTqsPwqqZR08u+f/+eCtyipTxOrpdRxUHoo89+8JQb3URI11e
g7ZSaKqUX7U/Fi2J2S3l7iSxJFad1vtp0MpY4o5vo80bO2UjM7hWVSzXJWhVN78d
IeysR2zvL6C2lk7BtX45+9drDXs2+ZsMDjX3jWVO364aM2b2MCTQfSGKf9XeV0VL
UgiD0BQm5xpNvBYdTri33s/E6A4dinik8Lu4lIwy2RjG5XbfyL66BcWvknbpDsth
COx2Q4Gu2DkwEjEBWcaQuGg0e1x/NcA5cwA5Wt7SYqkAAOIkXefBY4D4SqdlD71K
ve2lcUvBoz8wWwLiI9wAdMr/Zyrxym2QrW5rTsnh0uBhF56RFoC8gYhtdhEX/41V
QTbrNy2+fGR4HS2Big048HgeKMmAihOGmgoEeW+D+JnxfYduhZkWm/KhSKhCZt/A
yw3YdGJ/6LXeIjY0FfTXV9cANsyZgvobqc7IFn6EpLItY8df7S607KIMFiMRQrlr
YOACPiWENn5HvGwR7OkeP/fiChmtjsmsU2em4ha9SVqKMycJrhT4O/NQQVcX4LmE
FU4VxIeIziSzfLVxadI7xFvAMJdEU3EUorH6hpM+9A+/IHnR1CfsvAU/9m6Crjni
2N0eaXT/FYOJvJvMNb4zC5ujEQW2mL4p74JJvGbqsLROIK7Q6rxrolErycACr1J0
N9QJKFr2EqrWXemF+/EztEjHoS8YQIFxmMbV672tlgqPasd/BQ94THtwj3HgmYZg
2yRODSKwd1nTm33gtCUz6GKzU2eBlLdmeMShccPw6XdgIxSf326A5YVL+FkyCuHY
VxiRVZd4/JupmpZ2sAAr3k39ze8R4GFpFugb4WT9UYZd/ioh7aeDZG16CCgvk9rL
h3WwwWCfYIjOCGl7wZigD3qrIfMGdhisGwuqO2/HavG3d2drTwWyQNfdorthKi1t
+NwHDxnEcurkwODZ8yakg3dpac5d9ZMOECdUInPbiPd1bHGJDD5PF2n6r9RlQ5vt
iT2iKIf0MCoZU5pC5qE77NKio5XNBygIAp36g8OVH+8wXMnXFuxc1qOwuDv1kOA+
GN60w8pV0812CJnV2cuPSmvc5b4HkNymVKuFhZPn6OeZkIGyA2ZnmNteXWGVTUpy
r060NhSwOkORoZhMGf6vi2X2mv+Ep41xrYxpItfcbPQKAPVZ63oqcQMOSu3E+JMV
OtIdeYGsSqITycfp0Jhirpf1VDLs0z6D5ojt3tkC4a2IxDf5+QR1AemPhReK6ARv
i8hlDrHbZ07+/PUJjNZRI+pTQExCLjQc1aYayok6+SjOy2GN5noY2XqQSvuT8vKm
uNcqlYv8Qdfekqjz1Xxitt01dVaYqrdLlJkKITBYAohAdLy83GoD380Ls96JTtzA
BBSXqnWIPKVla8MG6b64kUj1hh2Yg3mFL+XPJ3ns0iTlqJD04hdQNS0AGDCB24gv
3sBD6Axv97dvmEtQAP8QUeFKUCQ9C7WP8oOo/Icv+tML0AFVl21YeuFXTz4EJVy4
6pZKO2rCA+g/GE2zGNWYAJhhm9EplB/UAfjdQBTSTMKItuc6x4g950ldCKNbGnNP
UUzcU0ixQ11A7+ytR/UTFNRyEXcHeS5jPCn0GdKpfrgbTU2j4nbz9/XuKyA5fc4H
sKg26XIIApR0ckwZc28IaWEqZZSe5SK1GrDeqovTf08toTxxDef+BWtuUeh1PK14
QZx2hTywrhFWdcVY3qxDk6DSRPkHfkwdTlR1Z5VpPasp7cjx4BhMrTIzbdpjC7Mw
8ZaGPT+vcEWXIFNQGUoGe2tyofUeOb8OGA/6J+pNo6iKNpHQarnnLsppebpYrCrd
wZ1NmpFaB56PXmAaP5f6q+ydGS/gpBU+MVk7v3yH6kEIgGDvtg98aEuP/IJVK7Oa
q6vmyDd497Ok5xrf1D9zm6kJsLmKQ/V9mCfXVFT/Nf/dspeiWuDxoKlDjjSIq4Qu
ZwvIuei1tdKPh6xJm+MUH8ifxN+bQvycZ72xuyrZATvTzKhes6+wmbjTpWulAZFc
RJT7VZOB3MEj7uhnKBWrmCH2kuMBuQ+RzowkyVFJ7Aj3uMkGKZ7DnOlD8G2V/10T
iiottHZZesWkE58KU0q+KZS4IHHI9Ppw7uSGlrdapUqjj0NhoEqIE2HzVESZV4XC
3Wv96FEbcNyAJkdBobOSOxb56XOA/vELnBSM6dMOQpV6fjasUMQOrdXcIl190NUR
gI5azANFtx1GK8fyOdEf4Qcb/B9khlxHlXRA+f5NkbJGiAnyH/TSo8qxtpFWUl50
VTCYkZxbDtlHzqhaj5oyVdt6QgO/w4JTkbCLznOiw1BLHEwuJoukfv4OwqY3HbnG
OwK3Ex4WGV/dDlVAgQ0IOQUDWsqScdYZA6of64F19AoZ5jnfdD5+AN0qfN0BfHY4
dJRnidMpBLmVMvv7wWkk7Dg1YHAR1binqELS8nELAfeTI/xtLqZRJiptFnUKv+GQ
lnt6eoIaZamzpn+fWv7vQVCYVbsS9/InYvHfhRYHKFVsEmSy83UM1yHuSD2GQDk9
OwTgkba0bXjPPzf+sCQVk6WFpwyu4hufViG6rQH3KQoirCHXCVKH/czuEyyuMdwn
re61zK8RalGEOm4r0lVci53QAqJHLYv75/43/xiebpvN5tYqScNltdkxOGVNNhsr
uVXWh1QzCt9LUqUkch476aDFZTVpX4K4Dl/D58mCE2qyVWYsnT/uXOTRqGD47zDe
zmsOJgZknhEHfh8IlXDAUj4yRkIMs8H+DEBLUwyuI3H2Y0Mzbr9LdYcFJds9u2nh
mT2HvaLCU+8k0A/RQV79nft7hjtaOhsFuh+7rA0BnxKcqMePw5e3FPFGhIimx/8O
snI7Wg1prJn4NrHmto2oIhtS9VxE9ezyvzCjr/7D0KmpoTmdtr8uAS22g4DzEgvJ
nN8/RyscmMuIfky0Y9C58ITOSRQcTIzTWdEKDb6pf+nBXXQRlmZr/9mE3GTL/goD
+2LfrgM41O8+EnwLvlQp/LsOqg8ORMX2i3NThQPHYrGoVU90FcXCMPH9piaVrw+a
vS78ZUhEh03NNDMMMNEITq6fVTiaMYW0QrtLfE8faPfAhIeT0tY82fEELGWbOnCc
PssRd8w2+8ImrAb17u4LPd0ct3F8tUkKqj7BuZtrDkhGzGowrmVXiMLq1JtuaaJR
6nbD+NeWjhg8PgxCs68XVi8gKT8Mlzxkv1XzPkM7GZ4nhloCVlkFJ+oV7JxQGWKP
+6HpUGCxOJt4cnsS7dx9W2gW56Any1FwRprWX6nN0l0mu0f8lRUblvOw3zMwEpTL
NVzVc5rIZZOTnrPIMqVEgaFQ3YZyBSY08zl5CGoZ/bXuo0G4dmxrriPN5BIfwXLv
4+KnA/1Z9ZkhNE93odNHK4a6YE7CoXM5ZzsxCju1bOEhbbpi5agLJbHNZ8PvrF1W
2IlyoTz1lIVDJ/nv4ogjNqKDsGpJbtSA61F6wG7xq7zO/RMECziXBdvgDmTZFDak
S7hSrvZDcSAAIq0xgx5fos6ieBKiWxEZoS10VQJJu17Sx89eQHplWoGnmza+NJ2y
N3BNjAlDahIFgp0VJez697oXinZcfqNUfdkr0LuyP6UqIQeY5jYiUsZjiP3gBNIP
kqWXDw2jPLK8feebYRLRX4glLgd/VxFz7edue+Ln4iMO2VaTWtR1b5+RsTHSwNwZ
2KicIbyMREAccjMi8y7yIC4KM+S0yjcywGX3UBPvgkiUeifg+edua3N0QVyoGdpZ
XBjUvdpQ967tkDT78OTSexscFnSzt5Jsj8laoP4m/C4gOAxkdbq8OTGJtpb5+Qvu
u+cHqxsjNAVyXWfW7Sgc5w53OThe33Y8+QS1lmdN+VnZJ4nOqyyj9yvwr6GKo/Zs
+0mzBmo9QLayVKttak1YnK4acIotIEBfGfR3J4cvjtwm9aZPhlzltFdaXZ9+2Qk2
CukgW9hb8xYlX/ban32D7kCWi9GlfQaDHBjmn1e/iu8lnllNmH03PAklrca0RAPZ
z61gI4dyPxZf0ogVoHkXaViKMo1hp4EueoBGHeG4IJ1fLXFe3bQ5R80NnCjpwNAc
S2b5uxwgk+0ogsGfKoS826lJbLVIlF4aV9WKFavMqLEdatoE9gYRrSouPl2ctsj2
udGVFCuzuqwbvNyIbLxX/DvJi+IuiF5u2yObpLHcn2bmQXuVLxsOlgk9QtXJM6Rh
35yqgE/LCIFLpkgvixUtUa7QMQ+Gyjhny/ITudgaGypa6NscF0YCJwONDjbPs2eT
4+s079YPI9e+AJBa6iT1yuaqyspq7oNDYc1xqw3/1l3f15R8E3F2m9aKkcnduENk
eFXOwZQnIb5bVkB0BODGcSmMFIzxsWErFGaaA8yZrNwQiUmvpiILqa9573R52T2/
PUe2CbQCl9WqcIrNPzAGtVYGgNPlBIOuGVi1hmPXG/Lp72kmlRqBuno4afQohZo8
gR8GxKKXKb0fQp1W0HT1m5SepV+ECn+/izBRrSZ3rKGr26WXc41ocntf6LS6NHyt
nL9lT0uIwJF9B1WrG0VZfLMaylJ8rvD9Gu2C8g8zWx/w1v+aTf9NZlqcpViD6vno
FgbbJwm5x7gOp1LGrQetesLdVz/bLcZ7sFity9cGBqrS4be7hACZESquzFz7dFTv
TX992ppa2SdS0v/56te/iKx0rRZ2NvpjxLO6lR7CkFlVdQgbP4vZOw/hnMjInxg/
evgGaRqmLpKOo3G/ii4am6jMUjLHLBhj4WNTLC5WNxOnKIsY1/zcZcC3yiUOuAmx
XmOoSV/SC+3/0rmerD71a9+p5EI7w98C+4Jdd/1EFFZJ7dgG54kVzZsi+QiDpjGk
PN1r11L8coRp5RjLBi3o6n/RGhF2jBfZMT51kAnBtQhXkEbSxnwz4j2sGMm2Uvi6
Pb0QLuWhu+RTiL5amYo220gNOK/QN0aqfwvJdPbmeQI3IHVZoNS6KxWOVDHzRG2g
Z/rvmD+afyoPQ9p3EejZY8lTU37KUatD1KF9pK5/RppLXNkO7GJOJz6QccVIUpMo
475Sd4f//pBq0HYCF0t2i29/iMNPDozyZEsJGpx0cGN4H1RF9YEuTtRJdVLTzGgR
qq0QuqFAE8hAKAR6F2oHqxw2wN53k0Udpe0pjML8FG5F4rXkf+6fJl50f9vAODSa
foSRaq5Sul24g0RaHBb8AOD2cpXgwEeNN0UE6+oF8QRvgpQA59/hsGRoLw9DCMO8
aLRAh+s0LYBNWQ7o8xDznJnkLMKvKxXhUj815fRJLawhQ67N4dbqjPt4VqFJAvcX
DMcPhrM7Pl6LjSutGpBmr2Yq8u4py7Jq9+c8auEXOdJTLILNUw8JRhABMAjJt0gD
bFl9nSuT82iypvfpiO6uray1k2ZWmxQE9UYXs9YEhP3ejgG/2L6AOhbOaqgk4VuW
tHwHKvKF62nVbjoMpdpfFSoMtLh7wFjiSxu/MMRBdeU6Db+hhqaJgb8qz7CjCOt6
VRXdcHMRTn+bUybdvnME2URCSPyM51cU5l8iYUWvQ1cipWkdHs7LdEkfIfPz7iKm
62R9y3miu4UlbjBRuqM25ocP1Me15YsBPSIrrhP3dFLGG5LWqqBP1YKGggiKXPfT
CkyFi5RSK4AFTML36Xb9v5aq43OW4c3Fb32J4Bwg25CK6z7ab2vCYtW0gmtxVtMd
yKrQvM2W8YNrg9mLuiMgU/h5g6Qw1te/U4dVZaHbCKL+5kkntbnPRvgS1z/dmaUS
hsEAqlR68i/9CWPjVIb6A0rnfCi6263UB7YiFVHSCYjJCp9dpYocG9OTzFwogkFX
KRilnOo4l2S/2idx/Rl4R4judZPjiDNTp0iC+iYk5fZJBmOWllT2dN6kEfLYw2Tx
epbqMUcxfjJNRgzdtcXuwpScRNU8iL4BImxQ+z+5JlTtVqPHhcfhc4ksD1uopeaA
28wsPjdcBZODo+XgzAH/sORpy+j/TOuenxgr+ELioO40KTW8maRlVhGUQ1cHdjRx
AJjRZSnnxLrS+pHAoQ8QdKrsV63KFSV/EewoO2vBFvowpAvpbvBWWY2joUBjv9fw
h79ruygwpvsayeFhXM8a2ZOh0VntvewnTh+jZqIu8DodKHS1ua4wR9+RuSxaIRTo
oSHi6Qr4kBsyabp0FtEjCFVmPIVpqVLMT5g2spSM8crNK5FC0nuVN5Zc5rrEG5DV
GfA0+c16jaiJtMFCrQQkpEDUogNMPTrxx0nlm7xdO8sjZBVEU+qvqrD1l00dNDGB
d1GMD3lHUdofxRdoWs/EIiZmIss/4CAvQOn0xKU8vkCm41HqN2FqKm4kRDNqTCGh
KH0xDlEg2KulCWhVz3oAm4/gc5vAe8EQHE7PEucWfgG3leXn2XnKtjM5E/twNUHW
6ZgHsVWcunUqRENf9Mq+lu+b37htcHWVRgSZ7B7VZq5DOv/UNpmq2kVXFfs/Y11T
qmUmwNzVd1OX8pjc2lZmz/0uaLVJIy2tjoYI0oxy0Uwto297498FYO7Ute0U88gP
7ZDnO8C2FOENxRasSTa0iqWovif//tZdXdU4ehUSPaRKbhDGnAAtKrGWr8bKEHZA
bUt+IQHd/sCdvBMVz9eKggCPdnegY20bbWID8BKUhBKXJrNsGfTJggK1AOTU9Ejv
1LHssgfcfdbptQvbH/TqcK3fVvECd8LpyC0rHlRjDCQMM687LFaNSSJoe2VY7fn+
+PDuxNhAS8+pXaAWhbBINrBES1WvNsqhRIhToipQr0DqW9JRRR+sVi6VlEmkGLl6
s4jWNi37KF8GJ68T8hnHhsjmZ2Y5zNvmlbmrL+valZoZoqhr/z6H1ViS7LDYLAsl
UO0fAi9Lwj85qWCFUzSBWAUfEe0XHyiBSoBLeAX3T7F/fL6SeTCHAg1X90vgki1s
3CoZIPsFradaT2yTvd2851e5QYGPc6nXP5XrXeT0aLQJ2uydcmlKA0JM12bG50ji
ThwCQRm/jaMQZ0XCHEaoypVMGqAeuOVGMDtJAIuSusQymjj9Djeu/QSTvaCWe9XS
1d/AM0tyKr7xpvsng72/kmLp2PydHx2KpCRDjKHcdKyGL+NT1rZcNvwJA8bv+IFZ
6LUu24NKmWXSeDsCsly0iSnbEDs5OLfwQtHPFhLBqM7A+Tq/apAnnjozRmGj+cUB
AKTZ1oR7yVNZclFyhXIqBSa1eL2Hy62pwdFW0OZnWjbxgZEgsVV5UWPR+BkHKlnl
QWHGXsO/tWXPnDH09WLY83DspQqYM5ETzDuH2nCeBXComxIKvX1WjE0gXqbmpn/c
7KSvoNwW81eYO1+qKgmace40sUZoIEqe0VLIUfAasFRMQh8IMdMmiomedqHXVv7T
utGUr9rW6GNvkNTvwKdGF2UXYuc8QX+obQnvlh1p9eE4HHF+4ZnWBKHKbKVkm0Ph
p7lgvZRR4K+Z96cA/o9GZPZXaJxg/hI8h9vpD3rUmG/RW+Ro2pwBAkNRQPrRkVXd
c5uyzJc9Dlz/Y6ZK8kAuBdgP9Ea4B4nQ/iforA7JsuWCqHKNOt3TpFR8tOxm/LfU
Mdl7nrgsfmmxiKQfNxJHh17aEC7toDxt1lxGUE8J9DlZQkxOF6RkaK4+gVBwyXIg
AVF2QBRy1hy0YITalot1pwLCGgJmRRBSJkkiCl1fq2/m8hWf9pcKC7fVLamsLwoB
q5+0ZAF4Hai3EWkxc2QYU1c3/7fhGHXr5wOslBMg7HiIZgwZQk5xF71mvGKLFfxq
Tdi88MRhkLW8BSj4ovFxB4p4gNQFqtINUoAWP9dsZFfRaqOaDNyYWvHFUnIFWpl7
l9DTeYlAvdD8TafiX4wKdPR4AF0eHcdc/WUIyPaXFwG72fa+N3LBwq6F14V5CWEJ
KkLc6H4xdUBUy5y2cSsTnipFlbuegeDoamQAqmB+EKgo493dAW4YT22CGYatGSJm
TH7lBP0QmU4gcZIcOU6ckcIdurkhgvUbaU2m9V82MGOw+aevpLIEGHJ1gmSe7RME
e6JYIpUYvP0gFIiCBZdoDxIIzVR1rqfATmfcrfI3BHVyohBI8lZVKQpjVzH3FeoQ
DoXRhnQi8G+kzGwkMGiRxN0GFYXwiLw6CXNVRHT3TMlTvAuFRdtIs3oFmOk6Zaul
Ul+c/3iIVQwJbt1ATmasHTFv38cOnOUEqBqdkjnSs8wjBvaxaZgFHJT685B0mpQ4
LkE5jGq1oW2p8huC4/wbLRL3gaZgtvD3/PpaLxH2wIVqIN51uef5n4kNTAjHc6fV
IEEFO/P5RcUD+z5bkDQ0fjZbPEg1BFBo2P8EFvapIVFYAYc4LncF61MpWg+SCbSD
ouyO+Xi/P1TEo+ruRzzvoBcUF9vZ9HRb/ARk98IJifCWrYvjcwgkq7o5klsgu1Hr
3Y9bza7QwJw7Un20dLDOTiB1MPen5iVoInquJKrIYoTcZKTwWk2SdBYX8Qy7Yegh
8AyQ0/iAkdLC4PGQXjnzDLlaig5GHtztueI1k5MhVvmOLqdcWQ6KzHnIcXsRfgfq
88YX8fZ+aBOLsVQWi9pbHlkBuo25AlsmTFm7pSobrFhnsdHpCS/GK1TLSIVqf9nw
B4y653cyI7bJtOORC1pr8Eojn+ajsvSn0cUb0f4NjL5FXJC6+i3wGZSsGp+zzBE0
3VT2ABkYblIqtDW6f3sJ/fAI71BM1CMj0mzNLWp/Njf2sJ9rdkIin9DkLQWWhZrG
0KN3fpnUXCLQw0tayh7OK5+TLI7H91NT7pzKXymeqkHI8M9NCT8uw9Z1bdLIyXdz
cTO245fZsrTHAPDDPqUlZW43GSrGExcviB8C2SQxPo+jAmqx2h2WpF04JdH0Ut1P
UanwxYDh1iltFuJQj/LPrkLuAz3009uNtZpOtUm3IqZfIUGOulQb47SFViJhvxEC
WzlxYK4e8ybtitxLnSTNjGOJtcYzfkVHQfVE4zmUUUYdqDygTL4R4Ps+qk6ME+WV
P6IarMFlx5Pc4agzwvifkr9O46gS5yEfLl4thSJMQpT/ovIBv7Oj8NGAY640srs3
sjegLDF4NLcrQArZRdcF3saJirSGLcv2UBEkvgEdImJQU6MnWqZvWg1V9afyZsuI
ovJ+VWQ639YXrymJD/qr8eNIl2eD6nucyVvRGSxbhMXva5HPq0VQxXc6JQ2R4v7J
rKUqf8tU8W5a0waePlAcgTBqXKv7PUyMUpBJvGWFJbWl0mqFjrykT/7GRTcD3ytj
xFpxQUABE1pCd0VCPqWw3OiQPojVURTtlhJDh4ZHHOPJwkSsb3iabPWPSRQf1mPO
651YiNg8e3Dd4uxF6j+HkoZzNACqa9bvC3mhbHz/g4yFuJ9LHYddEI4DCNaIFgI4
EY2X6n3Uvpojyo5Qq4OoMYjK7npvuHCTct8tc2oa1+Ki4/iWtSbMZN6mnnXAKIN9
1vjFe3u8q6eU2MqvYQ/9HdY+VIHjWFNu2lncocA+t6EnEX0CYIckyzWGFZZUWJFU
sSBWS5wqDS0jVbveRerCPz/vBDynw1JARFInDoohp3ChQto0iifPs6DYwiisarbm
yf7mDcEfkyHLArPOFh+ymBZwJ9LT79Tglf4cNYPVeEQGpa6Qaqw/A+TMQK0Ncz0C
45EPvX+ARCRUOv8a7Jh8GuGhT0mivSs8FC2FCUrMDdltt8UFtn0sz1JSxAPN9qeV
CT4U6M4Ku4NGLsNb1g5+pR79m+IYhFjr6jfh/EYL+KyMQ9FB2nnNYLfgIbsmZ6zD
zOlv6ZjpYiD180mxwH3TS2aFv0UHw8Bxrq3uk8EZ77TWxmzB/rasx4bxCn+QuIVQ
muQfQKvfwwoGk/iA93itaY3jqJxgNeWhmK4wbm9bkKumjQP1pZU1aoqrBnO9JOyJ
YQpgUCU0MhfGyyCJhwUF2qBXu5aJ/aFEjhIqqoVx0312Np+56rdtxGxa4W+NdnYF
Z+uAJba1LDKaIB/dCbGhNIwjaSAsbSUdcNWKGzy9guQz/DbNiNk+CPgxBep/RfRZ
bN3E6+xC1u4QG+pRdrma2PStKUVXlQBWAHw8GJhhPn56ApGHSxhh40mo9WWhzfD/
a9dFyg7ByuvA57RPR1Acq6Fu4y/F4UtAO193LuUIXe1WbC+RSrQXs08zc9KDp6C+
9OpE6ZDUklpMca/AQeU52KU1yTcWYv6txJm3huoCgbCymMtpiRI0FsMulm1I0muZ
5EqjYImdvlaJBeYYm0H2RM/ktbn2CK7eTxV+N7tQwAe4Po9oBidNqECnlyfwjohJ
btEc/LL7dxbvVCOxjydwnmVcJobPERUFbXsVAZ0/glY/Y12nBXjwkUsTgfREKkTR
/xLBSjidTNIT0YUPd1Z9US/uZ3ClVDvT9MS1gu6ZoBJ/jf0KruR3WUF2SYlXVxl6
qCFHvehQ3SfltvK6GMEoCif9cDb5fBwP5Mt9wirOBKyuG5kLjGJZ+MzVgdfkk0vn
qdCEwOddSZNY+JyNibxcf9fdXVxL1Phdpzej7Nspxgi2T4ofF8XOJd5W4wLVyxcN
wA44zFuLCCiv1AtPkIG3pa1xzzapjWFmV7fQox3h5JWI884okGgnCOgYdG3TWdzC
Uo+mM0SFZnKFBVMv9FpFPrhrzxIMMqf8BlYHzJYHL7khbUxlr2i2hrBClPK3J7aU
gEVnaRaEhpZ0KLIEigZj88Xqm3rq//OERSU3PWERVYSjvKmvBy78W/lD0PzT7ojI
Nj2DGhkreTBKk5MNFoyH7WGyqcR4uVhabK2e+crBGwbNLKLH9Th3j51Lrt9UwIaC
KyG/zhP3pKxk57Sn1bOa+0OfE62WxA5HoMHlNDfeHWZsRLwl+Kmvnae67kQ1BpyY
4/qM3Y+e+iu8TiMJx7AvWNdbMSyTHpHHWuGJtadiokmGzmqhX5Bsh0LlUPVA5LzO
LvA4VnfZXCbZVeFVSkgbGjOuQLeIu9RsM4G6n29s5ZCc1QngsilPGVzhpIqFfcYT
7NEPZvHE7XApjz/aFVpTtCGbY53EE3yJCvMEdQ8mP80bkcjQ7DmtyEqpXscUuNZB
KmXKdZSoCjUXdlSAA4KZXrh1cIlvXtklT2jZ3D9YaXgKWR6Ux2LU/e/WbLir8axc
mv+mZvSClrN+P2KkcDvMXUOT/H+6JVBTK4lGRdtGORyArdhuu5NtAKbr9rQV8Ufq
BGNo3ChMiDk5NKNO3NgFmxe7OSMCN3B5PkIIOj18XJSZ8srWlLJkqqhlVqWzEFSO
F7j3vg9H9wtoXmoVrviHaan3TFVHNfxLM5fyNcpjTkCekP7ay7+lcmXLsOgmvNi0
Zv1gxWgTaw9rNBOnyD6x1STNkSCNu2aiMXBW7VFTqI6mLYoSckA9nHn/ynlPzy7L
+4PPX2EEa5FFHwzST+bot6+MqojmmzHwx110HTzyUJMvtJzviSOyGqtb/Ccwl/F5
3yjMur6g7wMB8ES1rcpTbBwmszkJo7k6YRHYf2u7imglLHdRJvV3VTpuBybyPGMz
N+3PP5kcXYlz9NCGUh5HtYAJVBPLmBIx9XjYMSC0WZxYfUXgd+L4SWfYJfOodmM/
RqUw/5Tw8jc7ZZGBuKwuQAhVtqgfWmrzNolLhyJWepCN367C09EQhh6LLHazucWj
86TFyzvsYmxvz9aZY0e2oQB7ZRcgfsEj1xIotIYk3YaIFMdOahSj3n7xO0XE6I0L
Ehs6IeE/F3ZpF5vbJQmjs4FGM26DDIgTZ9kiQ3RrmNnRi/f1Au30jYQAmyYMsQOZ
RmlVJOdZsRbQTkkD+BYK+jLRp9BQ1+MyCa1A/S3ki84rh2fXs7KGTCB6B6v2CAqV
5koNh8RMa1lQCaySevBJoNgStLxOTJFytDPy1uVgCz0jqgG93K7s4j2pC2Kxl0vU
LNiOylhvlMH+ypdyHJS+Rg4b0xALB2qksf66HjTyWxDqlBfxQ/JqZsCGbV+T0MFC
uh7s89Et12eMZWCfK9ZxZZ3KqPKLY8IWDqSWjiG+BxH8uMQqd+ZwRGgd8xLlm2dG
R0s6TrVpEz5ERt/ciCFyWETObwlLXOWkCawkhYfnHMr9dia8IJK7St9l4YKGJoJg
ZK6tkhsMr2uENX3hL/ioZqe8C6oySY9QSKHfVZTuLXRtJSuJVrhte9ne2Tvtz6P6
/4e2S7Rs+AZ2Cdgc5dYPDAE4f0hp3Rm7Cs57tBWycZvDAxWVxuIBJyDiKvMDLzzm
GVfwLn/2/oJlA9R8uTJJ+DF4zBDeYwqauU8Vvwlx9kW+lEtE1qeeyt7krcZA2nvK
+5E0+XmumHuo+53RfeSj0aa8H1htcaS3lK0ajWa374cWIuOhCFEt435smFLcBDW6
fXoKaDZuw7kIX6zL16QHvzEGljULpvdgvHFqOBVMbSCghNX1LR2gKfmW670YrvyK
vhEWJU41+B/Hb7v8BbvqxKDs9h5LoMOOqsmwsiKcuSQPaTyn4eiXwPkBQRO3mbaF
Uoi8S5nsgc7rMRZ4lptrWXYrAp7c/QaEh0GrWHJifSrvFMk63d0fYZ++gUoz0Deg
ibBBG15ZYFcHKjr6XNy4gwyrI9FoS3xVcitkwySkyrq8FftgrumNJdCMFD7iTix6
p2Pe1uwEtVZ6mqO1Y3GeA0FKWMmZZJJjUJwRroAQQ7/TnlRD06y+j3m1Avi/PJMd
fMPQDbIMx5QElEy1w9WVv0ZKaSpctg+X99Sxv2/yVyHM6vAMnWNf8F7JxhEZzExL
fh6xzCLlwBeROHNpGtMJeTXlhY0d0UR9zhptng+q9U/KLTLzhLtemS9xff5STrHs
KXOLBwL5gkV6G8+5ReVsg0lXjoWiWOY9nosEJTtbPyo4kNHBHP4P25jT/bzGGHoL
s/BEwuLZ/jEaYoD/7mU/iGa194DYzwEymJ5cRZwwXaNI0TnoJKnw/IgIZnld461L
qs4v7LiWSRNZHztb33ujYvjyZIRlPNo3Ni+eklnPJ/DBiwkBSA4ynAAWqEquwJv9
r+DfkT1QHAP1YsUUr8GXqIufOIdrb/bHPQZsZQaWpOaLe0R9sjqAsvQmGwXsxhBB
odt345XMpDLsudSc02h1xB7SnVDYy3Rl7bI4+EZoj3mQYTNEhZ3P2PI0o44qBjFy
+v5ix68CQvDCr7qra1tjeWtRTZwj6DiyYiLQpwV+uYeMCnun1FMA5DiAGckuzYY+
3qvMfu0x8a1994PoTOGctA/+i8NuWasU6z1G0fEN9hxxR7iFCNqWJrjiegm0u2HB
rgfJw/+iZIVgbng/ejiOiECDphSDZmSvDA4uaNfFovi9+OiTogXpKqoIQvXLSf0Z
Ntwf+ZgQocPALXyJRJeHXnZyNKSSfD/5Pq5blNZHogy04b6BaGQWW1C6/oGZh7hZ
wXbE23IuzrsIU8YPV3Kmv9F5x6anr3Jm0euCqw0IB50q8lY92l+BGJ5/gxNQ3X/8
vlriMYYtztlSWPDZB+s6rNTp/IsWZOac5yAnKYmdIaTisPHO1CcP7RrlQ+8CHpQT
mie8P8S9iD/6GTQFZfoegUPKHhNjLJ+XkpurhNpirm48bdMePTSR+d3aONxW39/z
GqQE8XBic68ONBYuRWudIPIakZK++9JLvzxgv/4MefboNmAqFb1h9KWUXKqfhDRV
ZBgCZfRdFtnDCvy+KyGrNOXR4mBgUjn+t5sBl5yBbV3MptlFl9W3cYGteFa518QC
Ym6S7VHk2S8Xkr7JSBo4T0NM1tIijyDwP4sIHVr6CXxLC2Spa7Fd9I9z04wa0GYx
oExfL+daJrSjKh5vgaF4E4y9EbdG+r0QxwDKJGrcVtMPjQJiKINKuniG27JEHhKQ
+S8tTS+eR6HsLIaOU78fTessOvCrCz5ZlfTCU/8LYHBd02YyQfGyNTZHoVVWoLaG
aQSb3QlGdBD1gHkH5SEw2EjBwD/aBymcyNYWLtfIYm9IprPLZYMHuVISX2fudIPF
2QHGtnUwNfScRQpNWKZJqkzVw6HU9/ymrDdxiLGR9qAW6/7yZ4ANPXiZqorgbtIH
VmG235WGR1u9bTQ237B0cqK74XTT85ZvvntzlsUXjmO2IYVc3weY6TmwqrzMZJa5
DcTGbwYQZwZwBWvqiNd1bumRV1EJ8+eWlI/eQf68jYOk0gJB1kxHM0OIH5Dsi9NV
0er7KmFd++3Zd5Nad3F8YduSSLrKKKFurmcZmiWbC7eTw1BAatg1gaGdM6uMAXrM
qp2LapmHTl2DAOxowgb0XQYtt5zyO+1N8Zuvnx92eNR/rmfQs1Bk+EMH9BbKY0TC
oe1Hv9jI+lDGgABViRnCmAGz7v2wBSvXfxZtfaYOJ3YQOrnfvE4mWFCqSxTBqw16
UJtmp/5CuXNQruk7FyM1Sy6aaje1EjBGfKewjQIXlA6W5NLyGuRY0qlE3wR1bYic
YBiyNptQh+sbC4QltxTF7w3/wGB59N7d4WPagZMk1VR7LUl2FoO48udIG42dM3/4
UDFjhhJbWjjN3DUjW8RXKQZf7B6DY3tmIJIeZnjg4W+0Xohfan3imM7HIMKpKHOc
MnbLmthKu0hIcyJcSdJOMxTSDPrOOIeBGTotESRz4A5//I1crojIArHz4eP2MyRj
nrfZWhxiCxlRVYnNcktAkD3dLQfuc32Tw1kqSBNvOdE7qNJ0HMhEigrS5BsbidLo
9zmBcZ4S96wuRGwy/eFcFcfF6zBWpNO3zSc6J3/NkrSKo40xvKxdwofNxA/maeDl
pne4MeOYCp22cIRGJ9rMdKRbHjezC9ajGnoMEVSd2a/tqSc9OIU3Om1LdHJQEHMy
Fa2kGUtGAaZ5Y1hzw0DkDpfVS/C2QhNG0ABYq5pB0PsS8f7/N85mlLumIjuZIjbt
+3noNsuDuOevYfkvk6YN5bcTAbRYN4KWXYaqBxxuiztHoBlDpHE87rzn0N+NLZrX
kSqhwOdWG48QlUbfO3ZBXk64YUBBV3qscQpPqq/L6d3dGclS0nWIyz0hMLBO2/0+
OaHjruw8uxW2VckVumDRt1Grc5AY+2KqA/mUu0ez868lg/Ck9fKJK+9Ebb2Stg+H
wF1HafncYt0Oc16ghiI8+vlnwwCXdJAN4TLmNP0R2sx1QEaWY63s4WINN9/49T+P
/UfUDEtWu5osC6qdBhIGeBs4fdos6l0mZfZZNG4PMQlT+tXh1QL9dvIv8WtTL1Zi
/Vsm6MYzN9PewMFeJVkhWb5zPCLIBEXhCfpXc7PEv+CKWQoRyF50saL5lfmFPx2o
YKUl0hKKOiPJIBYgjej0Ac9jxY1XFeqGFH4p9db9dz6y/QZx+RW4YpRg4Zp1uBOs
PTp73BGbcKzIH2bQe7Gubwhj8ESRJKA6vdm18CQmmEp6eJWU+3jwntsUTiAwsG1N
vjfFGyr4LGuv5Bu6RsTRDc/Pe9WP2jhmKNAH0w7lBr+Co/yvti6E9cZmaL8vJ1kY
gjBjxsPE4Tfjd09ylpiSiax6D1Iotw627U5oXEMi/n6tuFQBjyFn5va4iIZC7cch
bfXtdgvHm440r3LfSIR4yWpSHqTV5WuFwXAeSuIR4iu8660VSJJqcU1Bk3EsD9el
dd1knvjY59ArsxcTyhg0J4gImEIa1KIdfA1Rr2iEDkBUq7meD7lyqobw+SIjrHxt
ey2/6lEF4VNWEe6ft2Dzwf49klPT7cb4gk/OXgTFLRQctC1rV3TbZIwKm/nzOW7p
omhlMO/D1+5SUNJjG65j/UfAWiuzlBW7R9KSZrdcL9+jDT3iCjFPBxeAvjde6C2R
vkIjjVziONMZGFMVFJgWiC5OiSeZ3n3i/5Sp6if9fDcsrUl6QJbOsCW612Jdm1GF
b51+gsxE4rYZFbwkjwQeELxEJz45uXSWNAe9HnHSkHmHCNrGB9JJdOylIo0996ca
TqhlsmmO6O7KvkO3ISAf4+2LCE0Ie6BVQBrlOu2FeI83MjboBjzSw9A9YKKeTuXp
86NMzTb1S5YvmSX63WfG/3QmJJBbr6Awqdi76llcxupm2d+1YToV5tHbcC5i3NJE
nsqHrP9sQ1VfOBQNa9nF6rN7aMKvttz902APIT80Z7ZRqzMSjZozcI0S5Tt9JSDf
6WEkC90L/Il4A977Rk900w4X7waG5vwwN4OCjuVi3uq6vchtJmnIBN73ODrC86cW
OEN5OHm6kTWCwo2TcG/19mUHKHovNOi9qdNTKuDymMX2797FCG4Wx3Lp2xZSmKBc
qab8pIevEEPRxjID7MCtGW7BqbVhyiEw1Hb4b1HjP+9Ql2lADr67hR+lyQs/8DMJ
XDiwPs5xCwVUxcc9RmN0S098nleXIpU17hX5FL1Yhwds2W6eVjTo89UWq1gN1dVs
LPjX3xb6O3jjy84+RnP5TC74kPKQvFa8iG6GHIpCIamyqrUrIYSs44Xk+tCOJP7c
wrmaroEPGwmxaC6yLclDJhuaacZYpR2mUyRy/74kjfMIyekChEPJerQFo8+jsym/
JBku/Ybe2An5DH3RXUhvCnihFuAQRlksLLqarBvapcJe9nI9QL7rIgPeztROG6yi
uncchY4/e7OTyx/JZHbOl1ojghSMx9Rq6xbOsHvK01d73z9umm04BNd1efKrxGNc
ZZkrobNhyeJkH8FDgCHtRgxREFPL2bUQmWKPP5CwFmcjGGKissarfaeUzjRpp/Ez
gdRbCnWZIOmAl/6nEiOQpf3O/PQcPCmzFH112NbW+tCMkWFXdiSpghxxGsOUI3II
pWoP2Ad8iXWMRLe9d7IsK8bmkehCiqdaEoqtCEw1HkVYHJCExfo6d/3Jq3r+Inan
kuBQ47cpqeG0+cWCaESsOko1iVx4qgiJHyUt9d9XsGQuXphqDDKEEODqqA+D8O1C
+7xfMNrXm/TYxkFbhI5TgFydUMkkKJjujU7ArAZ/54AutokE+Nu3N0XnK0Lhjy/9
s2AsY+VKOmQWhdS4H6mX2kLFy97wJQG5dGfKucY/cXK8vmaQd7ebry94gjq/uaz/
Jp7zDZldP9cN7Cyfs4I232fnuL4Ygd3s80qPrmdGzjzEDHsTaUDzyAZcTwPoytJg
TSdNPODGBFSEJMWhbWmyvhNInN/3VzVEhVZH5bGoMoy2gsGQp1nviMOSN/VmejJL
U/A/dC9rKX5hRqRr2A26CuUj6F5hoTpTP63Zxj2dvtrKiiIBbybr7os0f36duKIG
f18Y5z4iBiKxJA4tfruzpZVKFHOUCDiZyi3vGVs1NAuOwwoLitNDizUnRPY+qtOT
v4Wq2K/HPwgEkB7leWcghlCzfcfrWTZJJSh/FZsHIZKX0NBiAt3B3LB/tJdkuh1n
O2QwQipO8bEbPstzjIj9exXu644BDMS53eHkaT3ngynmxcD5W+VW3jqM3tc5h6y2
alc9n2KvRZ+ioRnAzIDfvQi2P4FfV4F0DWgP2UpKLl/2Xai64vr+MHE3rOks02k/
Uoh954uAWzp52+9Tf6yUm20mfdDyyLY59ML/TZdY6bbO/UNULX4GDGfSYcLF9nAN
XWy2k36idW8cUgub/xOtKuqW82GTCa8Xvudj2wzFsvPjb6N8Lx5NmzJK30RwonHB
w0voUfXPrAU8ZFx2c42OEetOA0GP0G/8JRsyUEURq/n8Y2o6sKg6z51pOe6lTfrE
MkOh8dA5BeM6Mzzb8RLs/Um3FlHUnxsiCP5vsN4tjORSWGTnoYoF5SxUbXAW66bs
UPcZMjvsCiZw+4g9Jrl/28+hinWpMwWNk0PBybdfp3DLC8SNht2A+00fL6d8MQoB
A5lzkuxAb15V3kuPhdUP02bQt7Ngg2mb5UYcFE1+C087GjZMzByFQig53/rM0TtK
sCMuiR24Px6DPW5lT9njg0X8K6DpsfePHo32WP5glsjhxFz8GMHFcoG5JpZAzntp
qmd41c4GF17boQ2FhyiRIzPUK9kq8l0aFiVtfs8H2rLFEP2nzSPEX3bzi/Lusury
jCidjsGqZkeTJDnIrSX/SAjw8Y9B0Sj/jP2k8/pmb+EnljPWrxbcH8PVcx17UW6i
A1KhsIhyaVwjsV4z0jvFe2V/Trlu1NJdDkMN25QMZo3It23DvClBt6qGq3U667Y3
SSVUT0/WaY6UPkq9ApAOIll9gAv3vLRuwAhTjq0nqzFFmSPvpiFR3TF0T7WJQOqt
xIysZmdelfNQjCB8OlWjgiQfONjx7dA1IbCleISMO5rh+G+QrlCov19b9QOPg34A
25L0V1fKjj7V3eiYZ+szwE946IwN0pVEb5ibdw6jlrt2UvilR4m2H6qbSryL7I7h
fGg8mJ19UDDmzwna3RTQLj5mjXd4AQjPhgi/4a4C1nni8yc71hvegcTfw07PFQEH
XQrlqkJ3bp9mHInMSbeJLIOmxs41hNKwlrKIZ8aJ778RCPrkb/bal15RnKurCz1y
HWnZK14LDEV81PE3qalYHfeuLEr3Dj+w+05M5nBRkIyWRVgnHaIYZVYx8djGHeX4
d/vok5T5G5gBjVPYyz/SJ4bkBhPhbhU5XSit99+ubEExILeZuszlfr45EJdt7fuH
Hd6WItAFgz6lhQ1wSL0gOifrO3VveAQxa01EgFfcKMhHhwQgNVXn0GbmcucLRNiG
EUx25fn0I1/VfdA7DOtMPExS6yaPNhp1r5usI91dxnV65IkSoXp3EoP0gYiSnbb6
Aj5Q/ACpqbyOw2/h1rsUkVfZ5WUkMulhs9g71dAMUvex/x9KSb0Jgaq3JQTqhnr7
0zbwIDC8+ykkzSs/WdXG4OBPv+NtvvpcFbUoMMT0PL3J2E8V6PLKkkrohfbLgJk/
boxYe1OW5GyqccRxz7O+8Fuhqvx08iFFcXzDmBWm247XscNNILHob+Ui7Mcn31mR
Ujy4/2rDqQIHHoEL81t7RpwAZT6912DGA/AcmKAMdFopDUCshPhSHHAm/W/fzCYZ
g1NN/QVz9aet+0ZoLiVHBu4G3W7RfrhnH0uctaxlS6qhn6bskceWa/UMA301A/yQ
CVmrwJ/gMsnXcWOHSouJzg9sKrquT2eVLfoa6CrVpN+JgxxzugtY7/8AcdSJ2L35
Iwe7HV6tT/aTY/R3xt54Hjd/yNJptmjc0lPYy95rRdWfC1sbgWuHXe2cuHQLDvUc
hiGcBhLV1DBFXhHvY02EXnrzgfJ8mYgnUKtUb3ZM0XooIwKrZdlvBnBWPF9+Uz7b
n9BTazQBbJZIR66co8ePeBmqUMZRg5hHa48wEE3ZrGLgdE66oJ/cMoim5GvYGIGq
HKI9Pud6WWp2zChyLgC/mBUfFdK7QCrX6GvJ+sCPTTdD485DThYjWajGUOWU2cAL
v+dNsOc8muiVDcX8RccWWHRQwR7q5JyZTD5IzJakHon+FgMDS0Hm8y4O5QQFsr54
rDbFDHJYZWBQ3ViWSPKppHgIHfgzh9rT/XMuLWpYyxCIPi0X7230KPbpdgMvrIVU
+UjiXWFlJB26nWIIPq5gwljZ7aJA8f9nuhXvGCzcdl9USt2jfylIXxifOPPZegGA
mRcV9fVBfj35kytOuBwRDrbkwTEDnDfE/bsfwRJYZGrSPHhrDCvcfCNiJlpu4n6s
5Fg3AZTSnOM5LKfqLqigaSlpN947SpX/Ff1wqZ9JZXV60XeJ8ofI7MOnK+r/ZjK6
mFP7wHrhrTE9FGBudIfIhrJ152o+Y1UeLl9Gn6znbTNcvf745fBQwSRsP+0I047l
UdYITrE1Sg4iMQ9kRWQxKy7t8X6oHvYronQCh6K5bVeaBC4sw5LNRZTzMUdge13z
HZ9dN1/DjK5G9dKWcktDc9rJSoe8HGHprePRQ1KJXhK+OUUon5ECqAf5niFgHmFU
+SGp0fGGyY0Bhibv16lcuCf0YAiqPUs9c8PPsqQMGzfXbE97evJpJtoeRWq7zyQ/
Ksa98kz/TByPj78VU2ikvXVV7y7NamKaROWs140zjlgof2ehen2hyhJqy+6vPESg
lwEDkwrYgVfxiqPjdPMDeGJY1Cb22/XegjzOOIgisudV61hub4FoVYUbxvJFvcjN
8A8cqd17L4/1PLw+PxKqNd4GhwlsoxhbPMqVynm+ZFHfFi71hngkDCvMsn73H5Zm
rUph5s+CvuRz2wefqBvJOAZRSopHVWm9BVWer2r9HebILp1j5sXD4Z/BugNLK0gf
FJh2KBOLuT+MAOfVdGm388iky0FBnjofuY0C5mXPXMBvderlUL204jQLJdNS22qL
2FwvpLYvcmfkXixITzg1daHqUmnjnfRJoqJGx3csCMY82X7grPE2rVHWi4OHiqjw
hVvRkwGb2ieDRgWZplVfSHNbaFNDqWWrMrW83sTg9cKP42sdopD0Hlbgb3mLpjMh
UFQFfeq27jBWYJzy9kH0+EfaJtsUCYnHQl2Uhs+DPyeSMamR1cPalmu8MFEAQVJN
/sby6bsvPeXmpCWAJyNbnbnEo/r+DQsBF3nsvBhW+Jz0hjpuhaCg0SUDBcCIlQlG
lt/TMlsLPON/fDZbYoYfUbtnTE0Crkcueh4nkBgjQ86094LYiOLTrX2gpVRHlfVn
YDain9tlRGpkZQ66jj5oS2Sgb+kfOSu5bfM3iMiNhYEfJYrfy0c1BIPIJ3nrul5Z
zxTbmCWj9N2LD/RG0slrheQCT/kanvl7shVnOclKtbqAjlx4+xCW/1V8FV7T978c
IyMvEh53mpSgAyfdgB59pLHXe00gZurEtlJYta55VkYbo63mmCgl/NTBhyUroF33
N81kNWvJub+6gZr6P8571H6k5D5AFVJa8Z9PPX4zPZBJC4fpaKja7c9s6qkddOyd
PE/Oi89JyNaQOyRbWFvVYepbqfhpPHKhMkzzPBKspL58IUnAarbJ9tgxE8LJhNzu
PJw0ZXH6GdwnU+0Wkuu3LvMIFFB1u2yzkA12WgpEzhlcFsvUGpLLuUB5TH/4rYlq
VyIEd2WTewGSPDs61tw3gG/y5H1RvsW4tw1AElXjBndbhr4fq4zei8TwoXKk5WY3
qh3QZwI1wJ5vd/NLmp4WPXdaII9BhmueLMDDeiZVpVUzQDv5pDaXdKM4OIjeZ8Ms
ISwv7x71BZILtz6fO9dk/ExvGytpMKZhQBs20QSuqYDTvyVcYVEVqCO/4nrZRvw9
HbUBgAkQAMgnbxtyDJiyf2NVNPcpGBL4eZNDRdKulYqiVqd1iazOTD0JydDxw5gT
biw1X75ZXqHLVUT4EaxBfle3ZSe3uQ2Fy+/dgw45r4iAVaY1TQJfqxB/Ee43615m
vC9apeJyJhaoHEn8g4YQ5hBYmBWuHSvKqQeIbU9nRDdzM2iUIYfLEydZt4FEdNrD
4uIR4C3S+T1KpH0e6HRkGu2JVUItIlET30vtFxwkkrBsSMObIQ9d7+IfzUjMY/EZ
ld3XANNab72ohn3Ul5hm4jm4FoU3ElpenpbMz/s0bwPfs/qaN9V8+A4zZIO/mejX
AoFfeD2+OlxpoWQRMN3u8Qb9h2UU9CzSh9QO2cy9RFb7Lr4Ha8L4wsgFc+Mvincl
0OuXvaou+W5mX3wIj8dISEVe/JbdyT6sM6wcGcI7SyR4hLrWKq2julPCWJZUU5ja
WUBVUpgyDKEGr0mEYY/RgBPk/l7dNEKclONZAkCw23mI3OOP/bYKP/sbtnuCo23x
OecYAwjekCl3V+tPYF+FeZpqMoKLRIF2VPVU839Avi9UVK5JwN8Ui+Dmags7IO+K
Xohnz7Cc6AOx+ZRjf7oyZZMmpiuWdCeENvc8h+wa5Y5GI7KLGfgQLvMjXCjpqi7V
BpgUHTooNDNY1bJOK8DSgFEZ6Okh0VAcEaGHtlsThCWVCMgbqDZ8Qx1DmWPYs14d
RaQmXj3tTVGwzXHxE4mOFt68zeHtXQRYbesoHdMbmxPOun+/B6PjLWhD0xdaNMh/
Y5gPsxbifc6TPYtytNE8gKeNjHEke0g+2n58IiJYPLWhr/4166s0OwclztaKvMjt
ZGekAi/TrrID13KEHFLZx842071Kid74ThCn0fQeSE31q8cO72T2FEptf9ScC6qX
HIkLC36PH4tcfnUOOpGDIhonkCRXPACg48iNhuY3W1k6RVLQ3lkdjCIe3qp0yRbw
QVNQuU0mCw/9QnM6+ysEjLGbnQlPGQqTD2WNkhh+Cfimd3QVu7OpNcYsoMIuVLGl
NEwgsHcbz3y7Hd7qNhbhuXNUkU3bh9GxKvd0Wp2yerwgzVtISi7p4f2w/vdsAamL
SasDGALDuVLovXgGXCuLCuFU6IEa+swuU2yh5tSNZ93rEsVDr0afGuoKL3TrU4nD
5wU7MHFFvocxnKGZVGTxmczHSwXjT6jLmH+17W0qzy3uqO3Z21pOnxf2nA+WHirb
eWzRjrRGLrHDWFbfhDYHU0fC3VDREI01wbmhKhxVt6tsDcXKS7+FhieHXLNSR8Q/
YSR6YwYNWeam+zsgDpuiW+9yzd+IdNEPzcpfrqynW5Afgyvvg+Ch7pA8MGiRiSti
IWh7PQiPWjtcYcV+Ig1alKDibjo1FSLEZas9ZsegrpOzsh5xw6TXkgSa3JLNw7BO
OfVuoLNWLlg9m7XF1ARrOIyoJgabFaB1PU3xFb/pII2n5LIeHks4y7QIi2M1OIso
5AvUV+6qmAzMnjfyiBC/QMYMk7styeUF2ysbaC4T9kX8WNHlrzaMEra2qIKFYdRY
mg+MX2m+rNjjd0kmqNLswa53s8PJ8hUSKSnz1qoAMId0/kJqzpH41zdOE/SYaVzl
Oivjm74RHID9rhdRlQqm6VuMERvKSMtzRxG25K9V3wlCgUPCPy8L87nrjKRwLHLS
DwVTb2YeLWZtz9aq/1tXcBtHZMyOnJi2lPyFfznvMBgMLSYbiMu6G9seq2agxdwD
4isqZTycFhkK9CUYktkMhkPa3/kLkN8shCqbMw3q1unw+iTo57LmG30exH8FllWa
L+7Q+vf99D694DfXAMEiUKiBYP0vOodWG5x1uqfcQAp/jLqbx5yr3rQC9DjrpbDS
YDYtI442e+CFyYe1RQ1T/Pha2C+Qohi8WIpZuARfDE4vppWUVetmk85vnrLtAqlc
TTjoe4q7B53qN15lYv5/SCroBmWO7S1ncI87Gu2s79koyC4uSDja3zr6TUYmWk8P
tpp+ZgHMw8SIeYunHXw9BVhBAAifl7ppfJkTfbPW7cfrkfADYh+J9KK+jo4xok65
5ByXc92HNKTL4G2DuHamBhxr1KWF5L1XgdnwzK/BXwMIywGW8t942NxtUM+kU4wH
wypzF/j3QHB9H/fOUCKDdXrRDUTKXe51ZOiHABFYbwlfJR8JJNbDoNUG7bGOd/Es
WJG4Q71Kb4NlyWp01ZOCINub9Nimfhbm7KLwBjPdTYe2ALBNA9B23y4QP7/b/tiQ
H7WC12u75RYEKAKWh3+jkyGVQIEG1xwRXMBPPkB9OitR71+Es0WEdJ9B9CVeWzs4
yMhyi3sPNu9bvS43fboMPoNlfPmfA4UcA1nWmx4t5sbikjagr6GOrT8syF+fIvcA
lavJCxcCE1SG/63vNqwcIzdrGYT57ALIe9pps0CJ5BYS8wsC+yNpSL159Jis/4Pa
NcVHIb0qCqn9bYfLB/IwGh8VBwkrjGbOFgNnAu7joYltauO+q3MXi5YMFgmCO/6q
adaJVQbLHi5EjdRqDspliMhyE63gvPmVCiTZizPG/lbDReGLyIkONN5TrXT0ry+Q
RM1AKkzTM+XlIROOq+s60ohpPMXllD9hASQgonJx4Yk9AE2AFV3PknTFXAI2ZaPZ
8hIK6PC770Q7q8cGBak2XmnZQkWRvINeSqOt/6EyU66umtemjzZoosnCnKi2WlUm
WQpFYj7fytcqtbgQSPt3jlTsu1/bOiQD+t1JAug8uBJ3qj6mfeVC+jrCZlmibJjQ
Uacm4OZeVDUbSSk5N+7LW7sLJ+FgInCxWYG7PWZDYD5X4y7gTFH8r81Qegav0yBl
luvh6Zul3ssT1tL9/eN8HAf1YKF+fJX5YrhROG0LXAgsUVl2fAg+6TNExc6o5t9e
bNuj88k+vXbucyn+w3HDQBdVp8pNMjqzDqSmsrsqjxAV/cpS2WCLatfic6oX0GQR
1fUHm5A9/DNFz4Y6qzwjuE9kTR1gtTC8asx04UN599HgI8DRPsfSLdQWqvTnFRki
49F+fvJzmzkbwCdRVJgkciZ7qKzapDiUnFhvcr4WqfYsSsO/gzqWoEQAHDMHBYGF
UfxDQJqKf1DOJSiXtl5ypbwnUFS6qhQZCEAdUiTER40Qqf/Ngx7uWyWWPxboAlwL
68en/Q3x1bOCh2mCFrxxPsD/BuHfBIob3wcq43H35YqZpvYoTbBTMKKYBSmTqb6J
QZayvaCiVFFqGs42mC9lhUBDboxRzPVLv+XRoVc7+1YWnnDujdz31WO2KY0/tsVe
cPweIpsCHCCZ57uZhi8m40U7cft6GmmkOU4YT5QhX0uVaP7SljQyTpevVjjvBu/D
7jwJNEIaCpVPmTHjNA+Qs44mBJZgWomjSYZbuRsRn64qPveoG9ERmAnIAVTyziM+
knNX/Gveh91pIJb+ACxeHK4Kko3RS+h7UwccQFd6BpMraPdbSbQ2laP5tboxHFCj
wNKhoVXotEBX8H8mGRqOq7iCo/396Hn2t+ZPsm4KpaPSkt3OLUHD2W8zCDZNL/Qy
W6MPRGXIGnK0V0XAhah59VLwkRAnw3Jn5F6O8G4dLoKyy5LzhRdSkYbQEtR/XTyS
8VfCPYxYI2ciZhsM4DqcqGS75M91+9kVapNxigSAJRrV31NFJ7YF7++NZS079zr4
Z8IQ/TbqEk1Hs2slGAV75s1VS9/wi+f16rsAH83OGvR2fIxfY3DGcIwH01HLNHw3
bCta/5HrDc2LN109HBRovZ/KEocDQ5OkYkxzjWv/KB8TMueUaRB1TUgVJwBaWbHG
SWOLmu+qWLhJOfGm8PorAeMa4STSrUAXWsq6HI5jVA6+g5HNF/LodYzib6Z+uARU
Z3kSl3nqlSvYZK5K5LzgZeaxizCLjSnbsUsTGA4s+Y5QHNfVxTV88VKxYmrPRMiT
BB9Q3KAqsgkGERYvdIGXFRWeYynqsVDbgc3r/nCZSMTGo93Y9BTBO60ICBjxGKEu
kpFAgtoKz/0X+YWDMRnIxg6QRFXvdj3Jg3b5mNbiEa4xrxjjvboACBkDsncr58ZE
SWBLSoK9kUnEaDuh1WkKVtEhtXeUsy+mrhVjkYR1Ccl70BH8kgBEtP7oJQ0WDzef
ZKMPuEcgBLhkxPsXzY6EORXFZntuv7laSn3zSDpE54lbpDpl1bPCUjfax7GcQZRF
u7qmIZNvot3xWbcA4tODUkfyx6clRME3sxTr+lf2jhYT4+EUW3PtLUE1WjntMBcA
2hA48OHqrlbodSP0W/4092/W1PvA25luCnMawA+/J6wDynftWdQJpu3R1erf6elg
pm7zESzq1ItAJdrsjtNdEO05eGVMdHf899QqY0+SaMqFBhje/qhmi3UiHWX3imkE
+m3UCeP4LBfp9s5lh9+0P09rFDi7eO+lfPUIrK1EQJGr53k3uwndjagPuF/n6N/S
l7ebiHi7b+G6IHP4abgLLwH56BSKUoEJRF1Qd2IMwjtAKu848E0MnZhlYrx+PDIc
0T03adryNIoERIeBLoG4yGJGl4xm++vVF40ePruVOfc/Nnaftm8KvTLcq9SbAwJJ
QVmF13066lLU1losIQcb0jdes6lAMROV6vXiwI3QPMdZxUdagODnY8SbR4VAOrLs
GcHwJ7AhFKZksa6pEWC/dNoZnSSbNziUnLwslgXlcDjT6zOtjKGWbMkbw9sUTU0R
C2KJ7rXBeQcud1VoZJQiTILq8QUPNoCfooKIpG7de3x8+IUWefCmk6umsgXKmVbL
N0+PBrcvFLsNVeurPCqYeILRuC/4qt5nNRNQ5uafgMXa5QVKDKXaYxQlj/4kSg9T
rF/38Lqb4tVKZEvZbIbbGSzBYSY7geAkssgf5TgnuE+ny5YqI/XdPRXFsYpMBbk3
mcnOX9KhEcdaQte94YhgP5NZAVzln5/AI0GynJCD3h2MOTKCo8NbpUtuge9wFgep
gokYYFkaC270OSxuEwCbxeB0uoGJV8dUPVtz5WAGKK1UmaEsagQAtgsnQEQjr//L
4PUFccKdBuDBAerUkX7zH1/yrgMuWS6rHIkS6BtVjvzmAICSTE+5iNxM7rVqpxhN
uM8qFKO2k0aai5diZi/+JViQMtedwHEw0AG5GBhRHXNkg378tROqjmmxhvkswTQJ
U8O25R7S3JIyKyrd+KKrOpfpEdGdyyNVjrXjlg4+VlrsxbaB+vT50jdaUDXttC+Z
JqrKPEBVo5cCYj3QYGl8/OaDiyPvNL7OUJe4kDFCDzUtx/bh5pT8UoLDdR+B5nFo
0GN9ETKxpEbQSvGUaM/OT/CogHOK9onm00Zi5gH+Trdn3DP9byvQOynTSbszKt6j
2VroHQ5dePjsBCZYOw/CCCKUkAL8Sjbhwfid8Q/L4RAC7Rl5qoKNY7NtTwV6cr1J
zSV6xK8In2JaD1P8LWE8mXFQZKIH6Pcw/GXCbiyo8kMfvkAHARQTu4vqICztA8mA
a33IYCGFVSgGtWmpKrr77bDiuu/X5rG4BoOamtxfdnk5SRo2rEJnyoXYQyN2FYHx
DAImQKiU70sHJo1TlxzyTLJ6JPexfVKQJW7ICsgpNgByz/oWOPKJjYsAaRp+zLJ8
FCJaDDCOsveOy4hp40wEnLmfzsQHBp2rfFsIi280n9Wzz07F/Pcq7oFzIRc0Z5bA
XU5MPWXVee+m51bRibhrohcAmIa4v/gkxWo4gDeJtoEXy+Sm2t5gWGBdKtL1NdPb
lYG0k7FlWPQqjmgz/aR5x96UBs1T5uuInVmJU1hC2AADnA3r5qgGXqOSRegCLm1p
n+EbOWu35UvOUshVpFyTMYM1Q/mmRe56yeoSKDjE8LibPFMrh8UlLD+6KTZEvubB
RKVWwIBcdk9k5Tbwi6CJLbLdLGuB31KPnoANKAuVgaxQuVN+KlIhiK/jSvssTGES
9rh7/9yTcl1NnR9EHf3ZOpcsHuN6w757mrSgPz6j0yTlvp6Lqj2BBndSPx577AGl
A1+pzg9hS66/qRdA+y5bQhy4vkt9e7YBdxKWLQ7qaiOsvbWeeV7N1fMt3/+PB4VD
jbpOW56N3ZY1EFBwjJHWXraVG0ynYCZY8y5+PrJt4rnW17ljN+Xw/l53wNcqG+v+
ly+RwdMXiJ8DuzVi5QEIu0OGqDC8eobrhhO0/hoQ9nHPm1G8lutUjdNaTRlrFxcF
YXInE0ZTG8wt9GeFzPvrFiYj1+2yiNxBvByzcpbE9GLsGDlLiVYIwq4nhdYv2CtY
uqBzP7cf7aeN6LUpU1SVoYma5gt9l1LAZVVzo5CS37dvAe4lY6GgSVTIe7kW+3a+
1dy762fAgxkWoX+SfnD2sHetDFXKXmGrlc0G63XPyBCshl2YcCIlrtKo/LJZGSl5
LchTu+ByvVppve9aNrLwifEN27T/Oyo3D9npaqV9L660IrijapfDrMC3PqKjircU
9oFC60xgWJeWCkTf0Vx5lx/viRaQMcu7TcDshCRz2U4ce0KoG2K4qLmqJIbIazww
aVlD87Z9H7f5vBWL+bf74waVIacBkoWxu3ayNu5aOYo9oU4+/nH37TRlcWMJyKRh
c4qaHiCiEmmLTyMPBFmBthxFCONgOwoUMHREXpwjXqhgDja60UifO0UG8VevxQ7h
6JD5lY5C/v6CGGOQoePS3OwLyFo7+HfQD82zNnUO4Zem2U0saKgvpsg9Ggs/km9o
pvwKpvKZvNGim+QJeD8WQ9bnjoyeABAFucSb8zNAJjTJPGGTYWmRVc1dxhntLoL4
8wtgpcktRcGmFcD2DrD2ivCDsgZahiMNJCeVofygGxxHIQyaPKPwpnMiveYlfS/h
EYF7nyojfquCtSyV9bXkDvQqa4rGvSUdhg8dcqM0yjuKqAFdtg8ExWRMtxB6VZPP
Z32+Smr55HQuaiIsoXAomX6svy2cNdW8+tEX+ydYomyzCd7u25ApaVvDs9drLBje
uLNzg2q2ooXdnIGx43H5+rOtuoT2WR3mut4xY6oCkzl+xbLxqaY2N4pFbchTEUQr
CshYf/K8WltprOajI6nS4aao35ux1Bv55Zxi3j2XxjgVERf7HbKmVnGXDFRFfcY6
t4xTaMJzK9YJ7YXJYsnKaeAfseWTsXhr6oZobXwUohe0XFCbL5Dco6JnQDxLp4Ft
dZGzUGCuBCBflab2UfPmKbFxOW8s8/Gl3TYsPFX+Cl4Ay0id70H+9X9Zf0DQhMtY
pdMIAjWhpBkzG/Pa+7lesb9DUa7DPZodMjKU+79zETqPYKizkWVHbfdZxMY8vfRv
CPZo07xxfLajPWeApH+7BLFMLRzArnKrR2wlW8zO/+tMqUAgnxHVTNnz/eD1UJYm
ZwP1BVI92ao4j1ktEQSetB+mtZEIomNisZwfPxXjS7vRBfcUuyueIp9HX00CesXi
45u9Qxfl6dgBSVMsdSXEixK9005U1kgTEEMvon+JA6AjdneOq5HqxUG2Ke7FKZqS
XHUoMHeabZQ7knJyNSPR5ztV/ZTE4pPp6Kc3P54rFu2ijfawVu0pAX5vAcAIQInq
0fCEAsdgV2Akn6CqmVNZFM3Rgx73Kxol9Ya64rprp27JOcVP8u++ar897Xp2Ylqb
g6sWQbWI2UmdjcalFRwwA+oLW3UhafciVuEAkcuZ6sTVIA93dtMvPbs3Vb2IXrRe
t1IQGM4xFy74bos3WvoSH8tTnJwg4lN4xLPU/7PetqiehXnjwB5qEkWfDJdkXp5Y
G2Znwd0pI0Qvt7f2bAXkt9OSNItxns+1Rtew0hqkcsHs6lMM2jMkbMOcExpp3daD
I52jPjDxV990AYm4JuA6nLDF6cwrGrnuyYbCq1ypwqJMzcUViDCUTo1kMGitmzqn
RExdyDX6UDhH8/EUzivueYqmymEJj8pSNb5G2lMsmeqFfkcLuJgzUqTe8htesHw3
yfwP1l/+144PHCOdlW34SOKs/S7heTj+snmL69m0GSWaDfFKB30RMWVaDIiGPfxy
H7oTVn0XJMm7xuGvJbzNqX1u4/rOcnUEpoXa8XbUiIXZ5ftVyK76i5iPQhyhEk9n
LcA1gC+LiFfgzzMTIdNH92ruzvIKKcd/hRlE7aMc8h3NbtAf3SUKmXmhWJTG+wBQ
Zli5vRfrq7epNX8IMp2mSCGHdTujIWz1XAM92BCX6TXMPPyZ2gC0PpKtqnRAyqgc
dWv8EBKOibezRaHi46nAvdZmHidTlzqkCeGCmmkt+7XcLWDP32hTQiJLurmUZ7X+
xvE0avzHdS1FoQdw6EWiKyqmm07g1W/RBPF9Yifj0P922JL+/9G4RuTHiHN6sZ5K
I+DIpPUjU0gkTsmm5Y0z7adhPJNUPljnRsq2lSCyyUoXuzGLGrTM4ajXe7Y+4IMP
RIrgO/Z7XgvjPCLi5rwOv+BxsQqlzWWo7YMOhU4EJfWW335Kt/ySE4jPSS1D6Ruz
wCxQ+o//pi2/0a/Zdv8TaS5F0/tpXLJi5c6fP8pjqu5lO9/5DbHQXxHnyYAtVAaF
WCId+3SPA4iUCjESJyD0t2rIS+Q69WZlZoOasenF9El6AaQkJWi4JQ3LnqPgeRDX
33tViu1V7AG3LBU9X2SJ5nzhEeiFaMpTrYMdOxGI9oaWF6AJUjfvg4T8qF16bo9f
rMxhEeCJsPUfSDoRIxmYxJEJXlfIbK12BvWaoPg/O4AOQXeOQAQt6dlGdc7gqeI8
jY7frkuRmzIp2MdaCFatdl/xprGJZUqTH3EXExyrWu9veF2x9+FAmdgvMF4FPKXY
XZq24MAj56Fzo1rbP6jUStJgoZZUiS3MKBEFw8llWuV1uhyKDMoiPdBpoh/Ug4Qg
BQ7eRHcXNSGSOQpFzZyI4UMz9RHMm4wbSiB5odv+TRaFRdyWWpcb92wVxySiWg6d
JGb7SXBF9MfyEk/L/i2i9JnFM6h0j5/rgMRUASsCG61GEBZmBIX57Y86DHsF6QHC
Kd9+CmPmBMZGGaOOKUi4H3dSKmmIjSfKL1QFpUYNZAbUarUZ30Fjt2KpsjPce+Pi
yE3rXU/hCGNxZ79Q4LaBj/q8lknKpZGzRt+R17TLhBAIHUjpkishL0KvgnzKMT3i
FI6UiYnBYBtCqsBaOWNtKk3frWB3CgXTTZrh8yAQ/ti43fXwN+NTcFGy1HvXO0vh
e8O0DDTDPrS/w+GmRLZnqcC2v2ZjoAtySZF7W9Z+tkNmBqEayB6qP8QCWmwt9DjP
0m0/efW5pyfS9RzbtTY89oJBwEYe92L3buyWOkdc+UN0PgMiv6MNBHCV50D6BEoZ
g2hq02LJwDC82OCpbc1vJ4YByPVSWE7oF9ACSMboP6OI4pQPblE408YXyNgUR0bD
RcxuxpIZ8H7OI8sGpz/QP3h8I7p1+5fAyWFlPapZviuyJ74rELySHvsTcwMsPGSV
UJozGRlPMNu7yyCL1j5xa9JlUemxSqts4G18nKdBTrR7pJWjUd+Fj+qWiXZ87znU
/956frnr7QX3DfvcJ/UImJAp7XIG79I54u9St+4NH/WjbzaWR7NTMWRU4uhfBhEC
/HerlbumDVanQFYKBxIASPavciza/ASzqa5+yPwdqM6HNuiDjtIZYXAJ9mRfzAPp
I/J3ubKSTAYL1CiPuybuj47lW/AYiPfCTvDftXmW+3QglDI2By8lxuT5FF7bda3x
xlcAYfszDc+nIsLW0Bc1/skPlF5aWqq/qEyCMbQkTqDI1RfLygxSEAxATJ3794rd
tQvrO/vF0MByYmRuDUgU+dyFqTL31kVI9XbzwqQGdzxHkHUWT2jRje2e9eoCHfR6
z2ous/B5pbRZ9tF76DcxJpPSwxZ3eI3LcGHkA4vPaQKMa3+X1utk2fTLRY6/zPYL
jvu5CDuOYVB8oIa+v2LlDXsQA3yHGmNzdPO8XZg1smLDClsoc6tCRCR9PfdbRbaH
uuSkWThiMxccmijSrZrge3GHnMiqgwAICQ+1jLZ9WshM3BeJlhz4Dqt0j4bSuR/Z
9ntx0BMGUcc6qDenfJDISGeOgVovw6u5aZxdstcgnvu9nhDAFUGSbdv7oS7zDt0A
5H/PCyoWFGXNmTivH89H/J+KYa5x9ajHAIYCnhcWayEl5BVBqnapIKRS33mR2E8V
qm6A0p/I352HYQ3JrIcTHr2PEQI1o4ocFjvFNSDZcNPs2H6D67rELIxYThiXz0Yu
pwK5rKdUAM7Mf3teTb6ylVJ/rwsrguHRfDPF7a0YH3yHOVsJBn8VmkyOLA+pGD7x
fPQCYfA+kySls7qeK/NzdqoPgApRMmbTOIpaKOOcdFFjtBJew0JL9QLdgFOjJS1E
RvWkZoF73Dx/57bm3kilnvGl6daE4DcsY8DLK9pp/fScC0PZM057ncIlOuV5jhzi
ICJ/+knIT5Y7KrFmKKaoaUBD6qNCIo6YfbOESEcJiA7EtP5TQx3PX9ksXO2hfvtF
cnObLN908G00g+AS7O4Tl6pktlHgHdtEmpzUlHWYHQqfL2R2Htsa9R/FGwgZs9hc
sdNMW5wLZUPsQhy8oLkZTKkRgtyzHlzg1RqC9End+tAnRlBCXbRsrFJm8G2Q4fiD
g7OmUVH7I7OnzgevXnp8fYT9IXyrKyZ4Vz0VZwZHebF7eJsdvRK+qJ2Lgv/0VGHW
X4crF3hUXeDZCKQo78H/mcmO1G1fifWXWu5icw1wd4tcwQct/Dec77vpGkMKjfOA
qrIK3moyCIr3mocg3rucmXrFPFHJ+sjVbUVW3afjwJBmkj0hQuUuVXrA85VBejtz
dRPlkcwS2gYB6oOoss473UPfgG94XaToZJICg2TDWrV5GQusc/Kq7cphHYIYBi1a
+QSvB7K7UaGEAcqqqfn1hPD4ZUkOEl5BFmQxsM2dmjhQmEzP979KeVWQ3yx6p1lK
BH2zfXW0RyMByjX1u+floSHsmBt0nCGlxs9x94w12Qs6TkB2TUrT+QZogmQB+H1r
EHoiKlNs81WHcsNpKJ7hywS32ZcpQsp+wXMgQ7vNkjrioOea3l7a6WOA1xipT6ly
a6uOU+UZ7zoNZhHtPaUk26K4LAGML7ZCndb55D1NmcVAxmjhTcmrj5pKx5C69j5M
Yoe1JyPiPwTHWHht1kAhSKy59EC71gvT9+qJh+jtf12FokU6f5ithQU7nEZLsv7/
aZxM2k7YKSFKF4qxItEnWyaF08cG0kkJN2A5D4tj+HioYbvWk57gE3T7FS27H7MQ
v4QLSrz5WH2+lNwaF6ahaBSW+cYytHT06Tf3aGpxJ3vfw79+2z3htX+7n19dbP7K
GDF1fCOkGIADrGuuYhMbB6mDygq39lBMsbvklIi4+AdakV8s5or9X6M9ihDPcL5l
04e+kj1sdlyLap1ZoDgzMuYGei7u/mZvrif2is86y3hkNmnLbAf8rkJrXbotCNVS
TMXEdT9q1TmpY+AW8H7BBybPuv7tE0rtDXAQzsw7YrTADy5SajdVJMXLnYmPLpXo
SD2KyKAQ9Ah+QtNlJPUkGjrQ6jU8Lrh4S8BIMAZ6q/N7+irL6YYe0Ep73g1lq0EB
sidMdvce1lQyHQ1vEAJBXdifFlL4I6Wu8EumiAagLUS8Sq7tI6AQAjZqIPZ1TZZw
dLRUIZHOHqqebY/LfnEP35J2gRUAAowg74zECeFEhfDek82Qr0NCa9vtTGcpbCoH
wlam65IOyZMkohWXI2+523MZJJ4F/XPHYCDpeEjFbDXVrfMEP5JvhHYVOc4qUX5Z
H+5ZNnJDUcV1cTrCw5HpVVfDW52qILk9uEB5WZFhz35NZuYluVuVmoGtBxZmmHoh
aqI8edomKtze+K2PRXotf7gGAMOkRMmxRvGBDLsCtB792b7sucznqNirr4byCg0+
SbmihY9PFCRg2CZkSTYgm+u6jo6c1u7+w4QKJckrRmaU7bP9ZcpyW0eOfPv50Jfr
peg5MiMt9FOLOg6O3R10DbgAprDaYlgNpXtfVSfPYsawsEb6qPvGbBQptoMkPq/9
nSeBiqkFmF7d+V8Pu/jrAoiRZduZHOKxcJ4Na6WPWtecQIZZYPZfWmdl4XMkJsIe
pSTFskVEw15nckxLPeaerXJacdm4XXGOHPK5MRQUw4StWIpQjEbf0pPGrTAnkJYB
7TZTtuNEBPoJ6V6Y9ZX22JVdK7ApWzsLytwpYCQi/qVRdRItAcBOQgNTt5hZvtj9
gfJDqNoR0/LKHTwkeqOqCwyRrVRgKNqbRmTgwD5eCVPhTZO1velr/W8WkC2deWqk
Hsmdnzlds54LoAjRkT/FR84rMSwLEbFLxizhqPedvjek0MioQFWDZ01Tpk+w5Gpd
Td5u1ZwUs7FT6pUuwlN4G6rzY9F2FMQMVqu/QBmaocXEC501gkYTOKhIIVhXVuub
hh1DJk4rhz01tNfichjhZTf7eb8AQW0mLApLKy8Z8XvIy61IIwY2itPqorZva84O
V/B7WXg9Vdg57VbOEcefO5Pm7EqgE9g+T4/ioIquQaz66iumTwOGLAL4R1dDTOPh
VYh9q2G5aPj6gK/MXZFW8BI0HkY8LMxSse7N5h8Pkyi1ar+gieuczbOX2Zisg2wS
D8CdpvtZS2AEvmu6e0dUybL6VBncHWypqClM4TgicD5SICbk07b4yRv/7205nRji
tYivOtlWp91Oe0vGmejxMsyN+fZl2cMxXMhdo6ahg39Zq+uSQrR60Hp64oOI7PoZ
wISio/AF+WSAz6u62lk1yIEG4LpXNw0MkynrvSHAJ46eVujkpD0XQuEtbBfjKlb/
Bn1i9gZ1y66TRN0Lk99qfbqA8Vmh+2Y05oKK7L3FOnkVk3thPkadhgkDr+5kyxsQ
xWj7UNcm0jYJxw/w3I1jkQJUbFIh1pzDYvGa2bK3RCU2QvQXAayt0VqQR1JzJ1sr
UPMvge75IkqRZEoUXZ6xHrDAhC8LeuRAWDjWmtZiolQHv1JivU+IVePS2N29s4Xv
+vMsW4IeWvNaWjfBHclSwl2G0NL5oeQ6/tm+26QBZVZFhqW3giPTXGijhC7ReGSg
wH0V/6VrW2oy+tlSpIv1na3eSb9jrXboTMjc7jsYJp1GyaqSUlq7IqBt8R1i/GHH
UtlfyHAInIKNxQ/OIxK2D3V791RDhgSoqXIp3Ym67GVwozUccK3O25p+JyHLRZ0d
KGa48cl6Y68N2P6oQfojsbx/J+kUf+nVFZSHEtmbNcoZJL67XUGtDCtrDDjquKHL
h9uGiZ596rMlmtNdlfXqnwas6IDr4dyKiJi4lMTU87mbCRMkGglZ7BCl/LRp98/W
3oMpkr4B/1xKPiWINLY3R2cyQlL+SKGk87jwRbpMswTnF16lCEK3jjIKEHvFDXHP
/tgMZE8647YUT3LfqKqlKeNDagM+iPkiXOupmyjnrpGBovQfdKZUD4uvxJDUZU+I
aSPMEOoAhdRYj6vqq4kBiMtQffLKMbK+byev3SnXVeMIy2LwP/9Jy1MsTp94f/yM
XA8vFn3Cx/SOVysEtzO0iYF0r1GZNBI8DkaBHM4BjhJuCgIcp+UGgKTKm1o+u1aw
djrwMW4A8PVCVZ8//lNtACwRJIUy0JAq1r8JrTQl4v1xuBXcjSOOCitJr22vEVns
OWt9AWe8KOjqx8If/0KP3RhW8SB1pZuiQ1aUPZmcYYxvuyDNgipRp8No6T1Mqthf
cRoz1DgImVkuf29nqX0eZZZ79PD6+J8MWFlCj/6yRx8AFbmCiK7JCdw6ikM0RGaW
stl6jlzHB21jGvMOazurjf+Tcxj3KtPevDzJa2BeWCrLZsNPHDSlbXACtnUEcjpt
DBUVALIXjHf3LjFzpkbseccowUP34/3rGI4qjqWl7z6qR7XD9AFo3Jqxt+GJiCLs
YUAcNPo+20YeHPJEXZpOvyCS8ieLNCjB/xQSYGdFdQR9uRtLxRyIBRJtPOU+Qffy
fmtl8Sq2Y3oYBcOjS8kmRwS8YUn3KuXueL4ZiOSTSueJClMZgfOXgGMFswPx/mJp
leqDnRHL8DLRPKHkiB9+KT4p8UJQrCcBIHHX48GsXXNinz1rAH6kpGaR99XaNiuL
3uDUdw4slX8s42XvUR8llBLnKEo58kF6aN1FplwO2aXH9dvCp7KZjhm+CFgPRqsi
I1cJ/3xtA2L7kkMB6IfdMGqCQ4WYWrCxtBkyY/kxZh8SvTSpLZCSZsEUoNQPUHV2
8W3MNLHiIxzHgDY76OejEVJBqzKvFVVkxokWy3N8kE4Y3VO3JEx7bUcUlxvNN7jR
wndZVr6RC0Oo8gt8FVVcaQktaJ3UmXvv06/4oihWAgwe3lqshNINIozbsNRr/sLV
ejtnOWNPvasYt82SNHW+sWUsNzT8DrEX1+9hF8KweG09bDX1+dLgm57caCxnFCTn
hU2MQ2+Lpz0yq++4ZPq02a/yMWkInqj60PCUya7lbsn6beErtk7rjznXfO7dlRU6
Rr/gwwRSlxIAVTMTaBzI9V5xSIp7q7YjOMrvUD77+xTpJ2c0UNbTogmUBY5XPgtt
JV2s5FniDaTEY4ldJKRp5dhIuFeNHzNW2Bs6GI4OMc1I2Qta5chbCBpstNBIgfFk
P1fKo9VaIml8mcLgeLoJL2rKgmjSlYoA7FqaqmDnzTQcToU6fY0yTZSdorv3XVgU
0gFbvJNPIPLiQFxMuDyixyEn6kCGxDXXscGjXYoEeMIZ35mBlkpJ2VQ1ZG6Q4RKf
oeJ3d2OgD1QWA1RxaJaUupU93CsIeqdKrqEp11Uvsao3x8vj3R6CtfxDiVEGcexd
JwRP4C1Ed9pqzOkZJ6eGqxuuTIL2XgZ7VDeNBFete5m3RavzSQ5qPJoVZ+JVWgyp
VKUtWOD40GUx+qrSGTkhT6C5+ScKwhtt4cIUwiVC1dApwgKryI/+Qv4X9KbTtzjN
GdsAYK0hF+W6NDgdllw9+sGm1dOTSQ9bSjZw+VOELPGAn1ww5Bjr+9VIx1OqBQQy
wcHdei1LxxA20TlfR2uFA1fTMj/Jtxu6+khJem4vS56VflmVH1s8F36M649HQ3g+
pnJvIrnJ/L6HJmab5WP1NwFyrxXIBaL1nBXZJQD3yACTdtpPE7yUrkgy7v1m89lq
ubH7YAY5eLwLRcS5YcpvgF9MHAhDFzEQBxIJyPdt+uoRSxjGHpVo88ko43xjEtRA
URUb8VawZkMVWluT04SiNdo1aB814d2EduXK77k5UYRNpX6VfiB2zexa+otNifKH
eEd1WSingTV//hh7+rQwT/owGlgvkVlGlMRY8d/tJ6rg9ba3yp7c7m0DZQ58GOxE
ddEoMGghqrEu90jWCF59bCJoBeVpo1sUo6/LzKivM2bdCRJq+6E1Pem30DvngoST
vpZSus9m5Z/m15UDn3tZFUe2oVubrWtCdIbxYVyu7B8tcx7+NETI4nDT+Dbd1VUt
TrSFsxzue9IteS5Z7lXT4pxGeUKpzVSQoiu5kgjLoMV762ZoDucDs0RfyS4aB73s
1+frGDSDZPpBz/uF9VLex3j64b2sow3qMHLlz95pkVJUvD+9CMByeE+/bLR82AYh
dA3dd/mLHqRUnxcy3SYwGuMpRBUm/xftEqMSlig5UCUG9Vqxo6CQhtjtkZJfeS5H
X16eZANnlcTdFVRV6wo120bpNwrR512Ga5h67maaxUo/zI4AGiTfFqQNyKaZlK/P
OEd0LHOoMnk/pMezuh50QsfJ51F867yhz51dw5XFb7pjINmRZ163X3MQTdCOoxZj
oITuffbYdZltlsTYpamB4rPu8Izh8rYBiGi82a2P1So2O9RULjTstPF2H2jfkEYt
nHxPSKFmV1cPjV47InneErwcFxZGwypN4iQR6df5ex14b2qJXL9xLXlEebsZEwkU
E5TLELklh7QEy3K4Fl2zmzoCNIN2ZIJvp+i2PcD2YO7tcWx7+R3sOl1MLIC/uG7e
8DiOLFQH8mNPRdWOCh1pk4pxd4rQNoe3icpin70OeMMq5wUkqi8x3BZ1Lc06m5ct
g8VCIl7Qg2Zp51pqGv45FQEpSlWp7sNRYRyRfWPoH1djIlIRV5zlWxn1ay73ArAG
r3xyV9j1hWYgrcnje+p1nsx95/jh4B8Mhb9fggUxiNagJuS7ndRxWuZgCenLeS1h
d+26g1AM8543KEk3LQoP7UYmXG2PmXGRoOPKAwEPXwahruAVvnUCHYJSseld9Nha
syYETv593LIaqqPLdYCegzvzY6G2SUjpWwQl0S92NCWUbLdXlBp+8X4h+wFMFHEB
HAxLZWcTBbzaeYB1rh2w65fpyKgF3cHxhegTPU+A4NzcZO4ng3rKNEvLGPuTHCUw
yuLi5zuHKhuAvZSV7drhf7CXXnKJn1rdjrvRl16fx9eft4dukeqNAOdpbGKP2KiT
4lLGWBQ6HQz1BGqkxSfQ8yN97vVU0xXGUJHkRJoQW2xnL/+JjRWXq6G8+Pmbh8cU
HGUidmO1M3//c75AOLO3I5llhd9zWGJpEe7wXIFpwUJDA6fI/aSUAGNUBk4/nMl0
j/oZYAPBgiEJy8iOFzxsIy+dSWfChSly51I7+xMMSipoAuXchBKwkdHmyXt+NV7B
LPrSzfjYo0VN+BoQmv9QF6kjloXgSA/QdzMO8I2HWeP/DY4HkDTAnEX3Exh6S2n2
ImUO02vbKuMzOQkjjadJ4NnTdLPISp76j+MyH4VApOsRVLeqd5f6FNQpiEFG/DTc
OVmiNuHez8r+g2AjIO7SQpfEd2XHM6iZi1xXzXuXy/T9rnB+48Wl3/jTxjwZJtC8
mE3mxVvRgeze/JsVqvDxa3GFmEdFs9UDtjklxGtNLO072EDlRkL1JF/XZpOuMZ2v
7LvetamVI/zDNBIhd93tkFXlx2LMHUYzOlqKHQCrUMerf4qn6/xD1woLbJT51g65
ma18KdShYEPaO/Ma0wczEC7VvoeM3w9jAb5bEkyDqg3Xav0JMAmoMFBAQQnT8+0F
dv1vv63b5/1mP/2OgWvKsU9Ts3IGTMyIH0x9Ntu0WNkzWB59Gry7i/GF5TLW9bbJ
wvLbMliaorcJ+In0tvgPhikYNBfX3fDJ/j3kvaR+OprqWkO1+VT4kXHHELAApkt6
Cuj8r214kDD9Ooty7qqY0UvZOat/W/+HpXkJivf2sTfy5FVCZYH8H/WAWzotm0Dq
mgMtcRauJj4k+S9Rj56CEAGbZjwZxoSYqt9P+ChoxrpYpzXZbrEN4jWt5lJPkAL1
zH1H2Murfqu7PRoHshw4xjfI3/FzGlIutVYMfcGCSGNv7anlZazsQ4dNTg6PWqGx
t9Dv1Pu7IrM0y6zChMkbso/B4G1WzlUXoZuvFCLmR6JhPQoVV94d/bVsxnZ2lPHA
KWSI0ESuN3v2aQzeffQ1OCYiNIh36VDQUS5sc+N/XzV73dDuh9+3Z3fiLyMcHVKb
+E/gp53yv29jNsuImlaQ0kGnhfTGEgGyRC5KVIHGH3fs0XgU+H+eMiVIrX5Xy0Xo
qiss+KWzWurkBy5T9WEmXBEgEo4aTJtwRn5s2CtRGYtR96oq3F4oQTTK10XOW74I
t6diKSsM6hoOOxd/SKsV9ka4Cm5/rOiNlkz+UNwdM3h1MAP3VZuqcRDWWwrK6POM
f6JLZValCGD0IQhns/mx+8B0siHHhtpItsn+8kBKiaV6eHVAIiB4sPVIpbCrjQDF
vBNhrrnhccJUcPazweqHVUH8N1JG50Hk3tHse49sfDI8EkHewu6QK7Ti6dNFIqMv
oWEnsl8ff3Gg+qXQasRtH3guM9YjNOhDoT7MPC9mO4lTP8FpAXte6O9q0X6o+Sd/
RIAqEe747zQJbDZAEJk5zOrLy4fo7KwjiphuuumhM9HKryfaXh27mdql7+SP9A1I
Npjxkxh9VOzDq2yHpldgF0+ftM5ZiB7ORfGVMyJTiRgM75UZrG+qMN+QAw3dx4Qv
N6IB9h5ulMuCMMsC8ltrsCZ4nDdSI2rYqg+PDcWgCM3S7rftunCHn1YOMQ6JiyV7
n6hT7FvYEObMLKRNdMfBDbDoPhIuSEh5+jTkxTE/IRYUHRmllpwvarXScHRn/JYz
mEXDB2HvfSWhT6T6iagy3GvynRhcLarLd8VuVDtM+YhhwcbDdWf3eCBc7XWfnzQD
bADje5zOHpHNafNohPDD9LEh35cAPExdp3hHLoXVOIkMF32X7eRGBDlZkS5aAaYE
QGum8SOC2pNsVHqAqkTDTzzC5d3XQbFRf6WghRylpjtm6LVhWnXUFno2yKdyn8uY
v9E+ihchG/MS29NFTY+8YxbNKx92xOGbSfTBXjSHbtFkS3JsxcSq+KlMyOAgbxdE
Mf2GARUBJADrGZy8m5zg9o0LZsf1zpPycZxRfJWZUYcqWXq2PQ7//bVnFei46KPd
+bHohvAP6nxH1UYiFVgVtZ/B4qFZsoKBnnxhsbomPMTdK71IYNBIJtnjM4iWkZfX
eDazq6MtLNoAYBEz2//DRmsP1gM85iUDANiezX9Thw0kizEUTyWUGELn2X/B4xq2
ZyRZr1vtZ33EiU7Ja2Xhgq0agEkaXJ18InWIpQ6ANeJkYlx4Ngv/AMp7VZYl+Ku+
N6IoRotpB947noknotVeo6tPoePqUedfF9yQrp4Me/boapqnS4HLFrGCNZk4CM20
pVF72ezhemjSSCxkCdDF4wbKBOZBFEOsqR6V1t5BjrgGGDP8M9qRyYT5slLg5bfk
AfHKHUOJSzd8hkUsO2YQdqhQ1qbCqhsd15FS66K0gqZ6apSQnb0DxcEpypAxbO0l
PrTmmL6Oe2xoZ438IE8Moi7FNOPhJ+UreCsbH1iAqjeZEJsKnlWSAK+GCTmy1h08
qVBBW5DZbpd2bPYRj/jgkW63oRmaAG9Xp6blZk3HFM2TI3HKi8JGlTdWSwLyMSqG
1jzFNmMFC8JNFjVOBNiMGzFkHbqI0lWEDZHjhjaBr1p/BHzot7nAIFjrB8ZjAGFJ
Bxn5OtU9jbm8+mv9MIkuiZRMNi5lIlqaB55W0Sq8umRBXVgyQi+WYtiLSNomxCN/
IFMxalqqUX1HKzWKf6xOpnQwB9kX/PfBIsU41C2xQI8b9VVTYp9WQMN2y3pkLe/h
gLFCBPalHxefKk11jKPQE3nqC6FSv0UUwhxq1Qk/vfN7xI5DayleuOhDx70a+rN5
kOaI/E5dUABFUILCMu3nJs2xpYRz2dNq9crTX8m0xXf8PJjfXoKnEfFx/R72zOz4
bTJM4zS8fWM832QvLPgSkQZieCsUsMysbzRXNQIZKLPmDnm7BCx0I7d+ON6M5WEO
7MKgOFyyK0zBgT9q+x+LjMYZpW/J9lRyHrtaSj3fhwuTbZJevhACAU6nXRMTKcft
bjfr2pWcSkoySt9d5+bEdTIn+DVQd156C7lVnsRgVcEbTwWtfKV20bIyHy65kLX1
tbNnrqnpdFK/GSL8Eb3N+EqGMp4M+sblAJXL47TSCizxrw7Q0BNxarUqo0g52ktM
PHrV7op9YQ/QghUvtmyEVmfRoeFMkU+NCrPKT7t80gw1Ey0IequW86OTKDeWgawz
XwIyZDP+VZS9StQdroOWjRoEndFdNw/Hpd2Sa6vevFll9Fz0E3JUoi524TOThUGQ
Qyyv7luMb42u35MyMdh2ITuKaK+azSLXbjORsWwRh+11CGuFKUR31vM03nnqC4p3
A2VKawCKR66MjAEX1l0og54/il7vLiyUEs9GWOFn8zmrkQhcGkahMEHjeddde3yK
vYe2B+yreRRrZbRKSvURGmb+IW6wtvH3DuAIgSmyN87LH8Zgjj8kVSsfYv7qbo6l
I637qMuAG0fyQXB5aUYK3e1XpCVZaZCSyexGksgHTq5ga2iebSK0x3acIeNL3U1i
9TpHE9ZXWvDfsGSqK7uC/qlErK2tfYCkOoCoWw5t8wFQ2PhvgBYDji7EOCN3xo+H
ZkfTnZDPCieAFK3DFgPIia4UNRSPu/oUsB1ccyTcIVdYny36NuIuKEnMvVtJDPsd
azjozw0U/kU3ehVYrOKJ4TRyfAiAlngdc6INk1kG5dceXdiqWgnVrrieTFZr54yj
Sl3O7IkizAt+fNU+vroQeQQ3reJW7dQ/s3VecXeBj/I5JXKUAecYIpebVoeFfpXg
lBT7p6Q20mDKAvCCN3GVnLJXe2IJ4KCLxHJmePsEunXEuNaQxTYG5HPu9BdJKLZ2

//pragma protect end_data_block
//pragma protect digest_block
k0nRDW/Jwb41iPpl+QeX8habl1Q=
//pragma protect end_digest_block
//pragma protect end_protected
