//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
cctQyjpw+LcwxsjMacAycC5E1hPFqubW4OWzq/ct3I4c6wuKCLxpq61e06RFq8VM
Xo1xjrrvLAQGb/5n8WPZJ8qm5VTm3Jla0hS6lqpKUdRwX4P8nLQkIjF+UA2Byu2i
J+j8ZzRdiaaOjDDbKfw20oz1WPC7PpELA7HnEs6nbkp+VCpuqGZOlg==
//pragma protect end_key_block
//pragma protect digest_block
8MLA92Sb5oqcTx/4oBpeqZr/LFE=
//pragma protect end_digest_block
//pragma protect data_block
wuTGFPqB4ROvmxPFcEcqu+BWTdSTuPt4yDJJOGw2Wew4a54K0Z3SjV+eF/HAUvrW
K6X99Vk+rp2RVm9RwTZ2U/aHaaDDJvzwPFgYChllBi6p78iSOnhERRWo7upLI2LE
1qXf9SQgZSND5PTmjFvFWpHWpPOvfK+fcGA3E/CcDs3xWDmW2w4SYj/7gFUoWUS6
DTAD6mmP6iQGDaUk1zzE7bTLeHG5nf67VfkXXI24tYDJsg8gi8mXt8Rh7lS6VsOu
3RcdxXqdQ3nt6LFcAd3aNXFeNYHgSKzF17IxUmWyfZF+EjvmSmYkYUDulmCuXkyE
u4sx70D552fVY5WsAKuqqJp1aoucCxmZHjb6QjT/kJ9PxfdQoQXUJzKPvWVJpMfd
MqI34TW3iG8vMwWhhHgp22dizY0/grPHHKVsYACEp3tINakWGt33Hky9bO8gW+Ln
Y2p6pR1wyOuyyYtP2vambIRt7KrsZG/xBPeSVKJMwZAQKxwOgFhA0DRqvdvC7g9g
t/r8v6E+EY5dO/U8LfeyLVQwDkCEmjIXs2iKLMwKsG9NQxhgg3nSlkAHjXY1oK9p
x+w/HnxIS64dHQpkFs6rNdfZCr/EfWvBl4ZTo6mx7dXo2wzMJhXxyef8n8Yms2vR
XEYW+8lEvD7LHUZyf6njThYYdwI/9mGMlhkEGCMG/gvG6JIJ3gpwCWuoHQIY6FaA
Ss1ZD7IHi7B9Si/vdlA/EmS9Cmnp4KEWwiNH9+UZktX2WtKqIaYmuL0lzSaYnKef
SPwh8AloIxqdVIiOU0r6M7ckhhxSV2wUu3o6jHj9L9D+5FD1RBUismo+V7nl5bKE
3qMHG/hAHcn0cSteGdpj1T7as/+8CQnpUDN/SvWyjVgtPqdG1tLejEbdFCbINA87
PFS8RC7mQflezBDJ5GayIVb+ye6vcacZwkyrfkxi+qoiJUm+GZaXfA0Y+f9aDGAk
zUfbvqrJta3aYr8XejgNA1OI389Unn9XOyuYijhj2ts7SOtVrUtJbRbFd6RsqMzO
x1fw0JBmj+an/LtwNdU197xswQAE3bQHPx1n75s5gKjCFmFOlWFvRkXRiHkhO8/z
Kd4tZJRJejmUwVuhExLkuodjh2Hg0kqus6CCNrx+Fr315C1OSYufjF1m/eVI8nle
y0BAJ+rw0LnXnl5oWAdobfqEU0g1DphKEpDsHB2GRG0JPGm6F61tmIjmiwWt4685
vz1CalWnX/UORchyaoFLit+YF8vyGE2cfvr86PsaMS6g7cyoapUXuiFYtnTswtG4
AkgEmcouoAZWJ/2KpjN9I2lxZLwryKRyZuoAlVNgylHNaPMWu2pWHou8XifhfyNV
8lKy2k0ejJJYdLW8muphRoMRmnYqfCDVh72kccqVb7h/wk1Z2XIf3coy/JXbfDvX
5BX3ktZU5mmR3CQhYhePZsA8S5ikqbcpCXgRjWG/vY2gO+buOfQr3TCQGgyUlJpC
9zLr+FG16Bur1dsmRf5H2gg4N4yM3nSHF7BytMBzglhoLW+yWOX16JFaRtGNswT+
ppGJ0b0CWE+w3jLYxV9biq9YlkV7MiigaTLtKe9Zk+1z72rXLvX0HR/46orGGBDJ
OBL+0t39MBQzbbOU0U/QauXFDMo8czfc7Y/NPMJCXwK9GQc3YKbXm+6L+15g+kX+
vcVbBVERuzTWYmTnLbT2Sel07Pu4P1u/WN/YtcfzYhqKBONLVYVFZPXg/Xcz2DPS
fQGmwwDo2d5lJh9a0PyhwBGbIAJZ73xqNDPUWc/JdAaT/+ZRuAfqLz/XspPNIJEj
SLD/8XaCem91rXg21rfO4/pOOAMoGgP5eVLg6jB7NgfNCN3vlYNcbvqv9J5HrQ7a
HWY5+IaECDhlkOirExAPIMjoPi2DQGBU70NCy8NaYai6Tt4O1xkv/peRVB9AadXS
emTN7MCj1LYBUYqWyXDsiTgzpjbU53tFtHnKqjXWuy9M43hwnE+e0NctRFRqB91L
1Qim0AbkWorFy7hnfL3Wi+YalJk38GASItGj/ZRtSHiSgoL8ZvfcX+iMlgSveD8p
0xZr6aa4HQNvhT5xiPrv0JGJopPxCdrgYm+qOvx+eUxt7boDMSZoAFAj4ACDdleZ
YkhVWvc6YUhenXLbYCLnvQ6U4UWG28EuQAAQFIBpqMgh+EsItIX0MQGlnfphVLNq
0QdiK00mVUINaOBwTCcqK+CZpG6+VYWlxtxDUWd/vEDSJ+EQC1Ecb+nmOZKerb72
3GCJW3R0sxCDDBu17f1THVi58DGpzAaw3bs0lTEN7cMMK52oAL7WlLmBGEpAN5BR
SiMMAP2McLnLw5Tsg8iwWxtJf20EFuy3hOvk0s8cW2vLlRnPOPENkt+A3eCzyjlf
LbtBALmIvf/s0CnydWioj6Cv1pUDsvrNfxhTERSC3wLmSJh76neAuh1KDwkPWMwV
Y7yppTQQy6SLuoh63lRUkB1Sxns8tGXbseXkNW30snpyKK4sdMDsjZvNLN3YfFvu
WPPURBjE03P/KeHVvmSPhf3AzKyyGWwlicp9NmQQT6+a7j2BSDjrt91HCyMdzQ+D
h/Abn91pB48XVfu63oM9+8qbHZ79GrSuUPRoX5ykMlWfYlHuAO3d3X05OM6mjFZt
H4s5zLQj69lxT3c4ZiS1a5f4S/Qizb8qHLdY/cj/BbhXMhf2zXaUbw23FyvJ5+w/
9Nj07h2w8ZzqlW0pA0WOMaoAqbO9DfT8kgXlj7zzC6t9DZ8vUkkZQj1C36bvfuej
FA4wOxSxDzQ6W5rVXncxGX1m7sQaFUSKK8u6jWUK6neo4g0K0Hnm8vLRkwo9OilG
NG4l9E74jtXSJwSQVG0Bo2Px+NIltAELMmcNCwGP3uykq/yXjcVrKNCBTy+NJmj1
ThUvBmJ48JcbJpUHeSSTcHETdXVyGlywOs4Nl6OEz/s5/ls4NHlUPgNdZdGOgFw2
MS+CaQL1HgwilOCO3p5gTleuK76A6HFKbW/JQ3IjKi3r1xTjpXSBC7yU15j88I+Q
VTAYMbrvsUk1f3sdfdqkSX9Oyh1VF8phbIoILGpCsADIelQNvmcOfWWK8PEyA6A9
08Iz7ueXLfvh0ux/IXehK9eDmsM5hYuJ3vtGOpmMpoKFM10GGYb0mXt71alSimLf
U4IyYR1XPkhfXCsrrvg79oMhXSV1uLUKiW6TSu5XdrjryhopJoKPMIFRtMZIXdwL
5Gd4gwZM1Uu1NDphhfpUXvrJ3WkKA9VlRm5qIwAbM5/Xuwz9wGAsFpLbcN7EkrmR
OsIaz5fIa4UneODkmjhLtilIcIJAJOhw20HlGjieATF+akVafHtuhA87pXHhPW/s
IPqRdK1dp3kXCxEtYpRAXGEYDwEd9IOEfxiPHnFaRdxXPC2+KiU1NwsnBhdbOviA
0NhU0SgxsSYuOWJOOt5dZYS5O/emMqaBOHNCWXpKjEkdFzhcg5ytWx/+iD1Wzyoj
ZhfRwdzHeZVvwIHOggZ4NtmQGDlXRBmkyZlrWiZWT9FWDf2b2K92FPDrczwC8+y3
j4c+WpKiqif41vgHaj6k4JnG3i2FMpC3H9Wb8ddW4LEgsavCeo3o7O8eOzMHuRJe
jagFDd5ule+zBMEch3R5jev6SicY/qNxYdkRfup401gsmp3en/Fvl/5luchpeZ0A
tzpvbgxn1MwvOoK9j4x9sfRyrstuUNyFUiGeoS8uxfLXHARzqu/bzJl/rU//znEo
HnzAe7MS1a6dAsz8fAczrn6mWfBRn3D48f/9jAvFbEbrpEGIhL3RlBdVxNMBXpRm
K6YQ54q//GvoO6+R8MuzLvsFTphOrDMjzElRuGQpvH4oKBs9+F2jOjvy3/JDCP5v
hxOqA3M8Q2nJly+pd1IfQRBuoLlToVih/NRLxsw7cyV5poWOfZgbnm57BNJhzorY
tvpleoOC2g/ra2Kii+UVh/nMsRmpaxJBeEp2LoHrA5sZyRDAhUNRCTe5N73BjBvU
RoQE1QitJc/zTqG9mc0xTihlO3ehqR9LFdmDBOxV2wTVKZWEsvYRdmVO0WJzg/ei
YtXtQlad30UaRullDFq983Sus/MNDmpXva7RrWHuvYq0BFBhDADWiOXO7ns7P+gN
JxQV3F7xgnF6k5YIN4rUMhUDOf+VfaGXfTbf6Zm3ycUlywJDMH7f9xAZht5QZ0kp
EYjKB/NTMOglR2oRsWOKSQrlO3taFXOjH5C+XZcJmbi4m6xxfgQNOFIlh4UHB70x
NrhePVPGcuX5psf+0hG42dxLDyUdZjeQYf3tiMRaS8ClGSRPsWyVEqG84ThXVvjM
knq//eWp/gm7pBC9iz9IRxzlewI6q9bVMZYk5dF2nNf0GyRsvw9TsLfA62+mkZcR
mSu3TgjTS+HThPObrAecEvPY+EG3kcWCC3/zkPzLMhcGymphDVDe3eSradj3hzuj
UxDTuLS9Uc/mDhMvp+d7iYbV8NhBi1yvluw02MELG4uqWDsFMcrExnFzNwam/rn0
JJjRJ9TFsSWNWqurpTRVL+s+gYYgFBaDodgcG9DPGOCj+7NoFQlEWJIGeTAMJOaX
nwaaeFHiRdm2NP8heGkNsKkiQ6dd9kxOQqryfCLhtH5LRB/4ORC90rmfNc2KAH6j
M+WZ9RqF5RmXDKmnf8JxV82aawtC6rEnf+9UQLNviUrK3zPiEuOsDbGuWX09p+Fd
RF21gvbde5iHvV37eFiCjMGUhCJk0xGDaPBVEKo4uOJ53yr17z+H+UL+vVW7l4Ep
XuXPapXmZQG2up4g6HJXjzwXvn/X6/XwzrMj8uZYAXRyaIuW0EUGy5XLZOaPE57H
kct+mpzlPhAGEpPPFR5b3TNTSTUdYOUYzF6oEMcrxm1GoM4enP+aM+LDopEYIqOg
cMA3tzm6BSCFb+QgA7XVSA4ss9LVmMO7EcgqcOy5FU9m3R1qipLIb+nGRLKyDTSj
yudqdLhOGkwS+807V2ttLADYLkKtod3R2r9LXrS5dQ/O3tcRtob7fBdZp8GWxUwg
E8g65zMQlAFLpIsNHI0RRUv2gBpmXsnbro0tGatsRcNzHkSL/Q6EZnmU2bozrV5Z
Q6rtXve6IDK/5eErnuLEALKF88Jb/Gpp03DHGyiDl80U370VaRPIO/zPps4VVzEm
dRlItebrOrszfKJhsptikEM9i/io9cwbSgBJy7+k13tanO6EvydoFawRXCCadGu1
XEeLcoZGQGp58yKKeCKftwsUoqnT6wcoE5ooU4VrrkZQpvOuugTyVM47zwVWWkAR
9oXquZlI7oqKGz3JpYp+2d8+x9u6zOlCHoimcwP6o+gdygfiKrwUpPkPjk0lrRRj
pZzA1IoxG3xBTcPwmwyKlRmKMrIgX4ycfG1DGJp4QxBR7pPJBNR67YF1f7NfBFMX
xvzhePVsuCJV+wU6Od1U0vtYDcuJ6CleBP5VFeDz3PmBO+szF5pzIz49jq5r6uDf
HQw50NqaFLZYvCF7qCAOz4NqrQoDi/hOTybt+nAKf/YLzDynlNmlH3EX4lzore9J
vfuCA05hQJArZvlUec+03yKbaU5TT060AtGhmnl4AvXxJ5hKnbXu5Sev/Id8UkbH
+fXoN3t38mgGB4vBZ/xkUvN5JmLlV8ErUlTyRy5jvytqQDeoaw5XsaX5dw9ZJE9o
kUHiZdaT/2h54VtfpDiXyR5fy8QLH47qzIux5J9KQ81XvGzWFJuvWcK0B9an++zO
RK5V7uEWnUS/hFnviycmLAE7vq1JZyUpsZOkSw8n+C8q50ZbU3LYdTrhn0tsmWqE
Km5Tx37wTQKyGG6haV6fxZWIZLicu1Bsup4d+buVMo9yt7SDAlNzPtRMtxFADEKz
od9if9Z5ugz0S13pIF1uZRzyqq8Rhb5ZJkKvosH3p6liJ71CSKPW/iPqtVmMcDCh
TsDm8I7qDLTmjfn75kFnBVTya1aOGu1A2ooMxFsk22c4N9FK8u4PEqbBxfWkimQU
yB9LzFhwOONTrTd7Zw3dt1tTayVpVctyDawjd+mF7bn7ITP+B2S/ldYZDgHv17gm
2rPDWLTpgzzH+dhad+LnmlnGy5opI9D2+q03/QexkHia7VkfnTi46QFMqaBtbRrG
tLAdOee1M+r2A01aqkdYTUiq5AXyw/hWDaQtK3MrspTE+vxf+WKtOctr2ePIsjaR
Uh85Q526wfpszIPY6fgCwc9wP+Nw2KpEvaESirC/0fmimhuZjkemfyNhLKzFLSOO
69McDpjJ+kG8TPaXwRIh4Yv0sxFO47ZzRml+bNsiNJv91QouihVwhNFFDYvVM0aX
SCJ28bhrJ+HYKYn+EfSRJazo/qbW/tVj1VSAXTT+7G7ileT2jHvMwNfUXE2qQUMA
z22HDcTXYwKlkaISJ8lAm/p703l4ptoHmdQW5Ey1ydpDdndEHuf0sanheZstDAmH
LB7PjJ4hcQEXp5bPnfyyQqIkhbw+h2f0fxilIt5uCC17OKK7VJilwsucywHlGe/q
wPCLdJK2Xjsl/LEkello1fapaJ98ELAqgtTezdLuDUt5xWOfh8OIyMUMROZ9JX7J
HlQEO2KOYaOwba5t1mGu+HGS952wv8ii2/VvsliteOUMat8/2Vz/hwmgI3If6fss
4wiN5bvVAtg7xe+qb5ZhcAHzdolytVuZ4hxcANbBBMsZ8cvZkixzzvxIXH4lvr+I
rwCxcfijuXeu1K6L5pROiCWUHBZLFi4TQ05+DmA45DPI6Y7l9Y3j0JyU1T1+UZJ/
EuBq7wtbn+dizGl4wczRxvQZtaAI6EvgfkwJgpP4E5yIIqcFGWjNbx3X42irWRpV
zQqt5s2dITrNN3sdJVMtPh3gDUC1UTMHu3koZrNQTpDhYcQqAz9A5xVBlpcNv9pQ
hjGG6gaA1FvsvTWFEMNJn0L+Zo9g/8R8lp1yr2D0eHNPfsXTzcGoZVT5SLeY0Tmp
E48ZBz9HOSWJ6UauRLTnxvaz3pJGyXk3R08OlryZDlHL+cV5ahAOwo8jSEEMuOl5
MJSNa34VJPFmZPAbimCQr/0Rks3phKSWJbo4VRugWtGkjFMnPNKE7OZH/wyE5OAT
MXwE0Ue4WytGRYuNw398c7YeD5IufPppDtqibPgQ0PkSlaV/fz0XktUPuH22tF/E
TNAQP6P7f4awgU9YIDfpfSBRmpopavSj3RRLNkUeD6nODZnQyQpEd6Zbg00gcOVU
wRK0lqNvbZB+z1OlhfR/WFt7k9sB85h0Zx9zmwOaYfsU1ehGbv4FXmAEDhaS/jOQ
e3CPcbpPZrE0QkE8l1qQums3q0sTyLC7qndpfPeR17M7Dlyu2Nkjs7IqlzUii+89
xPJqU9gMANNX3WHwnFoAehvGiefO0MN+QTz5VLdcUCk8GFvbtCJMUwdd5TOA3Yxn
GLaWzxbsXs4hqkt3+QOZ3BAyYZs5W7PifWZBVbeK9tuePcxRMh0XM94YNo5gbJjV
OgDU9AI4avBszguJ1mknFUwJsYVKOqD99NUmx/kuJ/f7lsKvTEVbyldT0mglw7XA
wgPUhnEQcu13AFoNx9bGYhbWjM3FX9hy+GFJxAD7GdsfdWtqhHAlqatC8yAf/EOC
BI+P7DvYw0tY5aCZB7TVek5VauXoeHmWwFk9trNgRH28ZBK39U6aydQ9C5irQd2t
Jtp+LbVku2CNUKznZibEBjmQY6ZnGdLhx8SEdLfHIeO7/q50aZbOLiDNq67n9Odt
imkN1hmGATwy0FKrKdl8aPQbcktf9QryxT7jHCirjxZpsibRdznQtK1T79OyiPva
HOaZIGh7SaSCDCcOHFVKjbgnakE7vMcnqiXPVKRP4+eyIc2Qvzcmc1Uh4L+GkYaf
+o6YPl0U2SI0TsI2EWYMHh7gXgJXeGXWXvOTNX/6AUBtaPqe0lzdMY0A8fJoozJd
Y6s5YW+/tr4l8XQWV0qCuIx1+YoK5GBNSbqeB902fy4Bv5P5pmb3YtJyv+v7spog
LTa/z6GvX99JSS7eYbAx7eMLNlHC3ZJGSl++zM90yYIH54bvuGRPWX2S7cEXGh5z
auuJ6k8wo7W9rgVC2z7HatnJX5K2wzWoVn9rLZwBFjTVEx7o7sCwXacCfjlT7Qkj
GIdvJRTWyvd0dXbF8pYCMkaju0ANVAv6xI6G12xngRwBtPz6KYrw0dQ4039OEOeu
0FXW4Y+9Ax69fV1nlJ7MHKaeSj4zit77oY2mm+tRYCxbH4DgJtpFLNrGHiSev/u6
zWxXuCTQragBRQg4htjAptbO9RLWa/pyXCNcd7Nzqa08PUtgnp7F7QBKeYGnHeKQ
Qbt5zyktm6kOK8zDQCcYYf0K/YWF9EIEALdE00x5Ax5Wc6WIb2Y2yhaS7L+Y2YF2
L/1LBNALlSLIPm+wF/cGNLEPSDCu9LBYcB/AmqRln3Sn8LY8Xu7NWM1xI3KG4nCZ
SYzNjyBTGLWJ+SptkNPGyxJyyrNGhusP6W6ekP7VPfb7Hs1IycobFZIUTPeQpBMp
jSGyd2tBpOFMHtscs8uYGfUg23OoXl9DiN7CwBNwGmE0d/1RBsiiHrLzbZr6infH
9a2oombW4zEDy5hRrWKEBprR2WhqstTN/RIQXxaDhUeQJkDOpeoSfP855azcymmR
f6JaP9BIp2w1XDRE6kPr3XCsF1tFwRp8UF3VhAfvuDf5MzVxqrGU3tU4piU9rCvY
aBGe347LnckFMF0cXd6r+MtJhPKJGJtfIBJbC3TFx7FXk2z0dHqApqlBXs0nu85z
anNnQz6EVkP5UqMBMJe0AdqprXGny0ICgjLHpy2AkuADYyZWB11dewM7ovIbiSQI
BIeY7ICFiJNh4LaBYvK+8UaJ7C7eGRlB84hcb0bOfRRC04j9QOoV860j4L+ecN4L
qD0ek++ZVpRhxTLHlaCNryR8owg4ojOv/oZbeHR7bncyrqPuyt66k2Rs02iTk0yP
owRtLWxCBjgv+BK40dAwYwZ0PYVG5cbaddia4pG5C2RYHgC6Egdb+jPqdwiADN71
j5K2PRmv7HqS10TLOuaNGbapItA6x5oo7LeXglJhlJxzv+n7HF3cBqr8xMYWgcba
nYG6GHaskouz8e41sAMxt0AniccT0xpoN/h0vkzPop0YaDt7Qc7VPV6m4Zc9UuUb
9q5N5ajJVi98bVLRjk+nlsycq/esjwOyx58A5OjAbjnDxBfd20AdDfb3rtVD99Le
2TTxKyUvo3TMNndGyeXEMfGDTjWdJrSVjFWUgERjHkAD7I2Oi7v8yD1TujRzW/uP
pc4ww6BBuPzr97mlBjLFy9x5CLCQtoExGOXNP1DpW3DD5RjsAPg1et6hDAtmqZ/Z
h5I1Y1D+5/CEnrLPEPGLfcshwMz1W38hGbkAcEQ1vcoUALMnUn0SZ5NyvThq22l2
rI6F7J+lx8eZ0q7EymwxgLSShwAi2C2IVE6wm4Xdu1f7nnSJ+3svNXFdg8HHlN80
tr6oc86DD0Kx+s1EOBf7dTdDE3wiScbwcy6t4X1SHe8xzBKJSsm4PK9pNwv9clpy
wKGsi20eBgXt8uzHVefWMocbLnT/fISi52kgGMQAWMLqgLgmQ1Of7d0uKPMZePGr
S2eYTxZWrrZCNeSCXGmmlNbJ5u/Zlt5MpznIq/wkurUmOa9Y3lCYzBKnKMV2LpLx
20PidA7l6nB+FkgJnLJumOiuhdAQovxC8FTM2Uz4KofXIA2nAtT65uaHRLv92flE
EPqJOPqyfKsUkTnbgGhhCzMW1UjqSY+Zcs9Tn84ke3dx4QrE6xRZfMMJR6m0z9KO
Kdu3fa0+02dB6OYHSyYCgac5xJ4DM8c/kmPsCnIdKkdMdy+MgIeeggxvzzl0oLYR
Gd9hoQzeohgsWk7tyMwg0BnBuBk9DSB1c1DhuMez8GDZiYiI4ubig1zT1qQkqOjV
fKkmylblGtuDgsMe57EmZsY0Jwc1sOpZle8PD+tkZuiVwBCh92CpFL8y2zWMRDY5
g8WqM1l2lUWfqrwb5rBXNwkO8GPg6NYZlA1ENkizpzKfLcM7/NZYbo3i7Na8IUcv
dkZ9dynHohEsrTcxq2yrzW5S8Tm5nMRVNU0u2El+oEMMEHw44+9I5kKreD0ShBHI
TagTHbUNQerxpBnpYUtGy4MhV2t8D6YDMIeY4WZpQZr6Jeyi+d9zNr16adwCnP0h
lLn7pxt/y4iQCfVgA+iSli578T72tmhNsQQ4xVzih9dYqFabx/FW3bPj2dD3K3pb
yGl7t4A5FPJsLHJadTSFqjuhsMt0xGCA05I/+TAFqGbFoVIRWiYF5tt3Wff20NG/
3uC38oCgowMWgukzNyniUeYeBWtgNM1coJKNmDG1ows2Qe/X/W2s1xc9gNVNxXSl
2+1af3hYQZ6Jl5teCMMn2TkPGAS9J+1X16efn8M0VQmisET/HD7u2cbyLgItJdCS
5yzI8bXkeU8MPf/cD4GVFJ2rnHMjXe2HtXm9nlUHp9XBUUljNOdTOS8ha6hB7faS
CR+VAh9VIlJMFfHU6DvW+1eJdP1WKk4y48l5eJgm5ON0Q1fc+MgQtvlpGk+lARcB
Z2NHk0JBCof6AGvaFjlWpy0wuC/jOTk7LO2tARSOCAvJZAhKWYGS5STo+JJ7aqWh
rHt4axzbD0g49+DD/vRCHbrPX2WosRWZ5qcpC/mxY/qfKbxlQA8oBgtQ/2TMGNkE
98Cx1VRr4UEniLMYlXFvFiqsVmoWq0w0e/Fx7rJAJdw4EMvk0uD4bBKMFRdTV2TH
HkN49ehL29MWtyVsTqgsoNypfqARw9s7hfRdodB2HcCCUJUvCvvI5TUbai7WQFSq
3k4N+h2R7fS9pi3PJ0MYegOXX9CKHLTQIX1enMhsSZpJy8chvlQxOa/qoQEyS1iU
881CkqhNihq0feL8+yneM/nvHqaiklr4ALVebHt4id2RGK2oQsMZBqpwv/v4lm41
Dgl8n54ixBPq5LUAwCFSUoSrcaSBLIRXcMlQIHEGllwJpTu/RW9R2RB4tO9VNJQc
Rtd73vnu8bhj6rOHDAD5hPXA8eY8QTb0kiflsNonAofzMS6LA+rjjmth6M9MIH+X
+63kCtg0fOlAWiX6qRg1j1w8kbUHzWjIHS11QvfKCIH3jw8xFfGE6ijXQnExaa6J
Ci/V3mngB7iHlDDVZjm8f47fvsCfRsOY75bNGnrMt/IpuwwPItJygHNjrsPv1Ogb
7ASSyJYJjV2wB4YHfPGpbSdi2yczm5Uuz+9yx1T19YuTy0JtEdHfGL9dXoEVfcGY
/DRrrQAMps1f5Kd4E2JVZXlZhEsLx/vgzd6o9Mm9iV8S1Ho2kEAvyjz2cpDppBvR
3PouumU9njwUnSRtuuQzajQwr/aik+fZk3pZSLpZf/M9sJNIxkctOElET6qd8Aa1
TyKu1vK2QcTPZ5SNC8xRTYbCMYDRUqDuutVfAlHcaJ18s8kr2fnQsaHqtfknnf1d
BlF7cRlVJLySNtFpIbQC0rHymmdKT6QMMOexODbny+WSh2PLBBnN8iwX+stV636V
aJpih2zfmzomaRhhpbU9lg/6a9kj1+IEv4Bv5gbekkWkJTDI82MW7pzfLdC7/nkF
G1P2pXY4fmzVzhdjZhjsVNXArSI+zn9nkiSLCwfK88qJkSPJnLPjOBfoGthwvuzV
KI1u2ASPiCd/qCKUJ84aP6yJEkqxZsg8UvUl6H9IKg9Zs561mxEI7u7dBxpN8JHc
6pLxw0uIlVVp16rWy9OD8HTQXNUvShbivJwPZ3yQWuaXKMwkaADqtSpBZBqr3Jto
yeHRd6o8j68QPAGqMCL4c5i6s7oUHt2AyI6McxDCFuk3fefkFFlWRhA3CRQGeVm8
0xXoSEWMnl1nBQvilcsEhfUd5e1yrvT2HYk3nIh0QvOed3TUoE9NIDQuEzL3zpS5
HwXH1+hY8zx74amEuqDQU5u71WAsvXIlVLnDRGK6NcjhjKSP3/cmH/JSa1woVKj6
feBW/VyJthhKdRZXtdjtkCLkujgavh6ijtJcjm0Qd8TCk77tx1URi2mOQa0C35Fj
MIEPJ2Vw4EbOIT1vYzGidZLKmM/lrnBeWhz4kqYvmb5bGvEiqUfjlYuLPdXOTnfD
+tkvJ7I5Om4oqXoPSMdfmez5w+sw5pS4pNFrDTLwo53fBRVvJ6J7HbfNMRLo0pCj
mPpC+b+qtXVO65T4Pf1QYCi5die0NZgRSLOzsgpAZoFltwRNlKWOk4uaEIjjsTAY
JrZZXKujE4UXnlLW4f9LbIvKNQMSLR52/BaEFLlz69+KjOWFjzFHmitR/gG6i4hi
CXkU/OEBRmWCliQ3BstxsrOsYFaTw3gfMdzC0hCzz5IucuPXE9t2pXLx2DDMkO7g
9HVY7sqb5LU9jJngALeN4j+5T61miLACa2t7RFH2k7X4hKoZl0YW4RL8pnNWwIRx
6y70ZMzMiC6yym/PlMLpN+BtDmpobg9IMwSTorAqUxsWcA+/gfn+i7wsA+krjcyX
pFDkdUZGdztJv/P8D+Rz8B5Mn/F3KvQBk6hJsNVjN1oX/R3KApoyheNJTokMKw8a
OcfZq06tdxLJFx+l63NfgwI+exmAg8w44f1Mo4kucndDIB3SF0/kDSdRBpTPMX0M
N9CmDnkVUTWw07JVhDYORZlUtD8PzGME6rERnWXIHkZUxA+hhRxw+kFFdwjtGrBe
vn5Wi/SDu08qgVEnADZG1mhCCl+tUaa+hS8kKyyhpfvtmbUnCQC/Pk3tv05mMNPv
/JDhe/ZERy824EPUfLK+wCDNg8fyE8X6E1Sm2obfGMtTWL5QBKzBZqdsWYitiK5j
G5cuNrZD9hsFGx/lUDilMxpJ06rA9eHurTn4Eqj5vPFj+0g6QPeYm1DrSWNHgBGh
neKfasUVP9jSmQKCnadLFDiSlLMtaxR7/+fiXojvuwiSih26jhOgRZ4115u0Ds2X
q5Glvt2lPI/yxLQQRBSJoK2HrRkfEN3nwllPC9CjQiwtYY+n81d6o0eT2sz6BWUL
ahBz6UXGGX3yCj4MXiqwqzJ5mQb+orr8iZcgF5+OY9defVl8aDj9dCp3RYuKdwxA
allYZof93w1/CTVh4VA0lFPBDd3VRBorfuYv5UgqjFD7AztYQzBuSSLV2JK2XivC
FY9Zhue+gRpfqIAVrL3xslOcIkLV/MXnM4as+k6N1LSCCkjzeuxJqchAq+vaRC3t
bGAEVSOqlGU9DL16grm1IyA/TEiIPD50yRIJCe79FWNHs/0ceY0kr4t+tbSXkNi0
l0S9j6vQMfZSnf8cu7ZF82VSdF/Z/G6OjRiya/JVfwwgiWNLJ9SwO0og7oakNt4Q
NYsnIc0pIrSET95ANR/fEDlQN6R9A4aztUSvdkoI2eBpFoSGMYo5SL2xRYq34omT
DN+W+h0y44K4Z//McmT69P3IsVburJSM0+idhLEtYj9dmTLrddPU0p+BaM6uw4DF
e2JYHDPsge49IpuzNHktmcUIp9eTLK/QUb9xleA6GI0Y27rzvsrsdZmK6vgqUwf4
AP3hicL7cIdLjWtNdQH2E+4nFTEuuAGOisgHjcVpovl28txFnLV2r8EAGilYRPgE
+RGCOEC0sppgddFnQnGQ6RE9RFsfnfF2MBGZQSxu370TlRb8aHLex95d0/nJuMXg
YSMOWCVijTx5eEdGChYvouN3Ntv53EwkhIurCxEcBcPgpqYCewOkMnkAzTo4tNlb
SKXlMdrVn0uQCxitOp/EmjIm9+ae9Soam0STmoI08XQI6cIqZLGLbwVv8ReBBrMO
wne8uug1EFENonRPTccCQMySmWKAhNSOoczDaUpFj2vD8f7d1iLbD+yRV7d/yrzq
BV2Eg0EPyHa1w9YmuBrSPNIf5Q5O27RBw6gVOTOsl8jaKh3W1DDT0ZlO48fOci5c
qN48mPp0vV5t+tGHplXJUCoPpRLmQ59vS9mvrXD4bz5ykzybT2Blsn1DEf9R12Qs
dK9qSpDrZIeDtk1wA0p6FbCARlcuRKtWoznzfKoXG6+K3rFwFV52t8qY2H2/8AuT
GJu7U1hS3FIMXjsMIUIzvpItdV13pihHrUqLomC9fYZ6+pKpBaLY6hcascDpH7VX
mpQ7TUfpHG2m1WGK+CliQO2BOwvMAa9GMyld/2kydMb5PSG/5SzoovDAZ4DBsKvh
e86Q3PMQu2oJWVNs2pYdY35HsS4HoCVbcY3cVmRvTqswGlO9SUIbl6O5owQnsdzE
kv3cyQiTQRbfpHhcdMi0wYelwGZwUF6kySqF2C930Kzu79v6VWIYk/saGXrUeUo/
HSm4vKMZ6ffNCcZ9q6pMgEYPi96nxiVg2tvSmbyEaeAdvk5LY3bz0/j7GNeVG6UY
djLptdUkOdyaBj6a464DTjkGmM12iAmeCl/COvtcZxrH8cXlTZkjR/a0bqdcMDt9
3cDqIXK8/Tq37rQ+feWTgOpWajtJGYbatIpnFHy50Gl5QoRAYeDqamszHD+6YV+k
j/eHmweRf7newnNkB0OHLUnmq/t/uTQPtZbclc4So/4dyQYvKHdvK0LpJAMe2TQJ
j2JqWsDk0SljguUdcR87FsjPC88EtULIq/CF8enyXit0Cr7/BLArKk6UEQrYhvZe
exyylRQ94+lsCJ+X6rZb3fOSYJ/DM63C7cn3J+ZEA3DQLcX6gcZ4MRKCYg1Mi/gF
XQXXYrYhJ69Tbkyv64eE0iM3yP3ONApyE0HUpj+QtcWZX0iuxyPjywTYMFAK0g8e
mv+SQ8iTeIqCoVj31/bwqC83qWCc1P0rz3FmiHkfiVX6gXiBgLnpv6fD7sInyf5Z
9tcKHNnwrY560WF7hXMEFuCEk+Jb1VaWuZvaoBMRrefza1D8Jklmce7uYMTuJGjq
gAU8/BE90XHgTSZj16a1pTCoEUydHV49Q4m+6FW6s/GC8SJU7OQZ3mnUCR62/C5h
4hXU5BiUPi/aC+5M5XAekZW3k8srB+NnOPDn4oV7j1cCLLmAYeNyCXO3T0bQ+yFg
WVnju+4pGDKLOoahkSdK+EZ0W/Nibxc6zudRjH/O3SACgTZASmXCmRDWGCiRHOx1
hry91OLrmkgy+EnOiDFDUprGFFuZKhbPS857YGLkuEruwaAU5/cSPAYSvmQ8oC7k
RYBHhNY1UkVlJVRRcNE7LIPI5rP0IufE6wJARgLcsuLqgl7FnTD40DRR6q9PbNC0
txmV7PWqUdS3yRrE15kfs0GjR8mhan2pwpYKLuia8RYHE2Vg1Tgghlllq+aU76WS
7VTXihXRoh+YqC80D/bFwH7XcUuPidhCU9e6x6UjkkfVYhgByvxkhDtxfhuQE5K7
QZkmQnWQKVk8dKpX2qXlMT8kZ9XreFN6uuCRe9PFryzc/Dha+faRd0+XnJFja8Ni
rRaQTUhr2JIbCZ41vKND58SdcBflWSoeoAxvPdJELDjqXX8hcIhiur2/J+otX/lS
jKLe3SBJD/yt73i7AmnoKtpNCKjnD9SSuS70g+JtMjDw29KyxsvcsTgGQ/oj2zLq
MUVVW7NXVLWwzPukKKwJb2NqAbYAKqdaJXshWJ2JGLuel03oFdsI/Eq4DEfwJ049
5VYx5KarGpb7xLzSNaNNJ2i7L2dE3oV3NJBNuJaIt04Ipg7UWENWm+l7SmkxgaTw
N6phBDWzZKERJFSdB9o99Mq7bkAxblBD8fsvhLNqGbW+F14EJO97GJRbK1oh/jE0
OKOPqq1Dp06XU0QkoFO6Ua6gVr1mlyN+2JuDyfapik1V8AR3Dh98U/7faaWQbrus
gEE0nZKiuelyhGYkVpTFI+LYb5Wku/ttThZFovBLu9z4/7IZE6US4R2+HTXeqvKv
UONiNFzL96OTiNCreqUIszqIvBADfNGgK8JyDm0eeY8X2MpjQ04MKvy42ktgnKo2
fgG1jHjCL++GacfrNH5vbaAT8aL+/adFYu2AC9FbSPNnMwipaVYtzD44AoQX9mU4
ZmV7OrzCjS6RMVae9IRhg2D+Moj+0XpFYJbVRoBQpqE/ByoJPPm1ku7ULFAQ2Toi
guIIbPip4pODeOCkRyPHpPUIIpPcZhjIfewkz33AAMnfPvd4DZy6wWTW42g45pwD
iqY5toJSYeSJdQGyrD109MrXJiZd1+6+aY6YllMX/5yxGVaoPJDA93sfZC0Oxhll
QnMFP7Ly7i6llQG6cfWnyaPgzz6+hhfkqD39p4zCUtKy7YffOgYkwLuL5KYE4Qup
GXB/bXX9K8Et1TuxLWRep6XMzR+lbN46T+X0UWl6QlpO+fayeVI1o3jqZC4LNBCu
ZImW0eSHSS5JAg7FU+U5LUByEHMH4QZz8dpVfjxuwx+Buxo8nm9Eu0zcCKNdAjtc
rVDyRK45D1q/VJqf5OoxpD9YhW37zfP9fb1/nlouZXNdJ7RKojuBpRoZJgZX8kQ8
Xr+hK+53RHt0aB4w4Yz7lr6WUdUS3PePltxX1/IZMfyVOng2wH3YOkLxix3zwLIv
3awBNHCt7zR47FfJq5EzazcQuoEt/pgSxhfwYUr49GvHIiW5NZ0gCmD7rUpGywP5
ER0Hmym7DhpcvhU07M2sGRfu4w3yaMCBdvth67V9OyKmX7Qc1nssrNXaPludFuvQ
beGHsZ0X5FtD6irkqjRYiSPOIy4ahclDxFE8IN9YhogVA+BOAT5kTLpSWAc2d+aX
E58lMtAPTqy+6IBi2etjtekFfstXPuYqwOPU6uHQgBoMK8FH2SC5XKG93lMMtZAe
fY7LgmXaV7dqcLGa+x38gvRnKJco5QcP/lNL/391s5szPgkO562/SF5VHmsdYp47
HQsI9R7M4nGGjdnIw+ZzXNpzmsEhj5zW+lHqtpk0Re9DicSCEzgbVaayAj7sMq7U
ZxTt9Y+wC9RYOgkUX5WQOzQdzkGjTK5PYxoHPDMjO1/XJu8UTs8BUZDfZnIeu9m4
Niqfpj++/Xiaq4kCcYCF2gBT2Q0WCnpWCJl/4nNSV5lKGViSOZUU5Mof0l5RD2DD
pebaAZVCEJ8nXRyCbgQccIXPAXBazBzBEALU5GcsU/2qjHY8DgVBqyrR733QlOJA
QnK0XbMuA0pjbhlWWo6tsTRb4FH6ifFO/4+IAfR/RSsEJcoWz+Z9sGsiu4alIwsl
iSKahTPArks4RaI1HfRAJoJu9vo43bErP4bUmYONRee9UFtKUPpeEYj1UxrW3avu
LEt0u+iyAqvGR7TDaRk3iXEfEEhtj3YDAWVLcA6il47ZDEEk3739nEshJUaxSiy9
3MaCZspb2S1d6ULLfY3u0PSqt3rt3GaIwXqJF7TH6PelRqoqeo4OhAUNAyGW4jGa
HwLjB61flE9jXxBF8r2Lb+EmalvRtVc0OEQPNqNZpq0rnOHyIBu8QdddlvHyBp5p
1SpsnWOC5NpB+9V5jBvh4CirKhxWSHL93N824SIJVMJ5MRUOSaVs9L1vmYklQRVG
VNDlHEREIUb4OzyKrEGXE9bm4PKSnv0Ip39Bs3ggwLNSYgdIQTXzYr1TeRPPPKbP
+ed8zENUT7VCzx52Y6IRUkAmDJtytz7ckUmH2dpGLWMvpTraJOcv/nsvckdLtFdW
DuT997HSBv87m5coWhOLySQo9zMKnjtlID4ahbrRgCktBoiajHKaT/5DzgwGDJ9F
rxkv76dm49qpVZwEgD2YjTrEzdujeB40kVj1pqc2J0xRZTluxI8SwLZkXLZU+adL
jJkpQ7f91P50/pvcKABjciDsHy0zn9gxHowiY9IK7M4Oq9fePvgxULC2s4bQf0xF
t5mAuTFgZ67AUpkEs05VfNQZSlB7gbNBWj0N/Ylbs8e1TRq2B7sY7skBzKk9xQpt
sIzsCKGrsd17Bhkc3P4Wj2dDU76LYJwPELXd6M3JRheiuopCTc8akySRPZpikzOd
7sXSArJQ05w/FcTdvSQ0kwd7lYGjcjuKgHk3g+wl10WafpcW0TRczE89Gx/kzFWm
vYb0N8G8O5JLdBqYN4kKoPDg88iOU5/YXAPxh4eR7zZlbPEoO4208PlUa3gkhFxi
jk0y5rNHD9UTNAhpxTedOzPj28ebbW4m/DXt/KJ4lY8zafk1Lf9CP490VA3suMGa
PG8LV5nizKETkOnordhTcRU5sOTgDPVtdwAzsLKWSjuPbGdXxVxchm/GgWlankmn
nIgZaZB1h+e76vJuCqauYtv5eQfivjCWoDcG/dcvWIWASWxD4EqO6HDmFfhTo071
2mG16XsrB6HtGBStuaVNBa3CODmr6Tx3q72nsZFZHMicgqQ2NN2lnzhYGanLrudV
CJKgndhTH9LOBfj3wBraW9lbNxJHPyvZ2RnoEGkjSx9wEODCNKio1qyrLYspQi2v
XZCH9rlBpBufBilgPKneEBB0Rla1+pdrjRuPQH90Bwwmv+mQl5dInCEFmMW+hFzg
/ZQQ22BQQqjLHV4/xD5DHmAd+ycrvFLKfT9S6gO/nCPKAYAE381CRzpatIjpT9vY
R+NLQG3DotJT/Kk3e9R8GTlCwHN8PpfNZxMYJmcTqQiP4594sCvsPTpwUt2uN1HP
L90hBiiIWLMYKX3L7CK8MAM19JzsX9K15iXZDaqEPaBbuOLquQV+WOj4+0EJd1m8
quOZVOT3X8PJPG3CRmd7TfkjmmnVjHJP+pb6bVFkyATo0tiFYT68egPCeTKzY1Pp
zo/ETJw5O/65aNB6ciTq6WaLRaHveFjvMW87Ut5XlfeNETupUp90LUm2DwM3Pylo
JoVR9q+kiFjoND4+xrGPdgcHoVWxJKN5nn3k6AHnyoxFi/bjz2BvEIV9GfjDjgO8
qP07HscP31sxDHEVjUIvFZ2jDVf5TAQwt+pr20vGfZBvD87n+nGyLO+6HJtd/lQy
1vFG6G0Ftfy/vd/TgThfNvno2FTxzSFGpR+uCIu55qcATuJqT/dajBy1WE6qaI4I
F2X6KTZcJCP5OURhRqZ4LSbT0ogsPEBNrywPtvr46Urbf/icl6I2ppoG6Y0Q34rB
sed+3xDvc9gnz5Jvyc2YHs6ZzYUB/qffS5OEKq7ii2H7WUaLCJY1axrmrYxwl9w5
bYdziNhl6t9AbGDLOYOdoY7AuXJP4R0kghzNp1Xmq10ZLhJiaROmJ5I7CBM7Ycuo
RMJ14YWkZpl9dvrAMTw2/l+/G0l9irK5O3BPbIeSi+TW5nG3Bx7+5jXjP6fq3Zyj
qYW3L9xl/gJ42DPdW/fXJ41P3N+lMQWmxhUj//S/Ci4KM0RzxLbYcZVQH5+Uliwf
gKKAZ04cHzUkjHy/8McsuEjddf95AhxTDzM3C2LqSLV/vndTBkW+C4yVMZizjclk
7K6zR3qHq8ciZ7w5HEfmlGQBNdILMgtyq6uFtDVZdRjiyHUSD77TrsKIE3rGxuqV
Yo5ydeQWiQmIuaw9LXhVkNhPhf5UY8mlcHliKz4zYl/Cc0DG245FwVw8Yi9IWPke
KafwzaXsWdnuqzr9OwiBgOXmSPQlisPigo/O0rB0q6yVuUeVJzUZeu8FcHBaPsaC
EbIvajekhWVQ+6B6jjuRyj19zCaUMQJQ3rCdlmJ9IDdtovlUsqiSphoNblmB+bbh
NCk7aZlgQ5B2KJwKkjE2p3o+mnV83he+e5qRs+yQHh7v/m8mbut7yAQHNbOUdt5N
y4hYkAq+9a6L71zndlU1zc9M6YO1PsF3rFr4t9OZCiDpNOYnSBexYH7w5xjAQGHT
1irkGRO2mc9I4bUckBCx7diQsAYfZv6wlA1ucs1yMxVhn9tn2UdT0L5uyowpI15n
YRALRP/yNrHQ52flz6h6szw+leHjQNvHiEDZz1YH7SGKcbQ2h3+uhr2FDNZztapD
I6bKXlmwI6uv7zCwJ6F/I3fWRZ44dPI/REHyyKGWJPWht1wCHk41HP+OwlBZJVXk
4+h9t1uxi5kdTAEgDxncs/n2PPPjIJ2nze3Z6wg5UO/A9iowViHs/DfAooYjXUeT
NsQUsP9p+0QgxjdBUK2Sr8PfbG7PBtzMjauJY87msvPnU2Tkeav/JpRyF97SqA1/
v+y5f+AlX6om1zhGZSG0KiToNkdD4bA/M3uFNoBpCTfzYcg+xM85pJKJWTUfQ+gA
5c3PvQJvl/GT1G890+M5flg3vks3Ij4f/5K6yFidvv6L6hSMm2Cm+WvdYFfbGvnP
pUpzBTUGdsMYpy1zLtyL74rhusUQ+J8fYbDZ+LjJLSHslnc0hCsEkUsTJyp/vIoY
8X1iY5arIxlpg++K6RI4743SwTY3lshXhAMndTqx+LOUCUwa0qzfF25YQMTmSFPd
YdoHFCRAyAqulep+pVbCxl9Hq5Mbta4HtBq+R6rojF32VpDXuywEpEbpgbRC/ekK
eBkSg/9CikneFw7ucQl2KJTlSolRYuz0n9F+iSTCz+uOFFIQaqTsbUZm8h/DyLyd
467mR6PuBts6GrzMQaq4n5iZsoDU0ND7rIx4Tx+xVaENvImpp2/XbYNacempZZGo
RsQ5zJtCpsu3Qr/XIaKJNtrImYIjl+m8UkMmgBKQ9IB9p8hlMgIKcQAMeq2rUD9T
A8oCnfhZD8O2/X971/f5yjvQoLzOKIvqLLZ7NNucOGODrhhRda/L80IVHnf7u+yS
R9+zAmGaheLxIygn/Lh8t4xxxjtE/fc4yWVh1WZFu9PmsTqy5ESmMppwFvke7WtW
XzKIhT0VUjnwB6NiNiJ0/9svYUfVCzKCz1qAwXufH89mGWyKgM5OruDf/FDdA2hs
/QM2tJcIy3ZU3dhnzt3pbIMJvMVgz+7ah745BZPrYvZB21JhQk1ZvtGzjdRZiRW1
ux9QSLXr76DSIvdmhwzggHflqHAskF6nmiKn9bZyq4lr/GHxqm9O4MwyxCk1zFQ8
0v9Cp+CM6ySqc97KBsD0Iv2qC3IKNehSCTrOH1t43QitzSNSu1WzJWkHm+VBjNkg
bHVkHZq1fKQI9HYPhzkw96rFFtfGC8rBjlRbHJpjeaHo9X0x79Sg4RSu4XQikvHI
lkc6xjAogRxnGT93qiJNZbtPkwIpcRsPnWTiF3x1dsQUa4qyxY/lBaPJULuae/Cg
vy5XNFfBXdCjisQO06wuN1hvDXnBih4M32S5g5vojJVACv177INs4sljRCU7n26V
nRLOmq3Wr8UbyE5aCaiGum28xYlJv0S+nM7j1xcmdwCD1ESL6Tg9fS0g5rWzPhGI
4c1pushbhNzn/rAnEaIq0G4JtZsQ2m6OZJEh/pUsGRuxsntSzIhPGx4JXqITvuUT
Yz4uwqWAmMqpBmi4jiKxXxPMhdFInaHWqdU5PaXWdiV04XqBtDAshkMv2rndRo6S
VgBrgdqCJLvBhlgIfx+Nw9dry6FlAekZ2BEj348ziEKESwbCD/+gK3swoBvyorov
7yXOMkRJT+uW2xytBu15yxT593h94U2FhpUY2FRa7RsyEOWDsRMS2GsZ3CL2dpBw
IULq8JmsE7a6Z7D3NcN6kCn+UraDsWCLXzED422M7vXF+KucGqOqPwP/hW9T+QKR
ivFhFwNLk0+1FVPLKEqLmBsLBNO7us2fFDy7yysqERoKmZby5/0wSBUUfw7fm6vy
J+hN1+yI/842ilA7sJ7eHidUOg2EgjnLXhu5DV63y94odMVXbEHKyIgAF/v1KK0l
PXZwcgUbiYbkuVfU7HkCtzt/pvLyehEGX+2q4mivV7j8FPadepfsWp0T1Gn/tATn
LfYnuajydhdWbuI+YgHFe8+zAWgUx+chE5GRHzLZG7R6yb+tZdi+4WqgewaboaeH
mIhRO+f8RJAPUjk7VOEqCSK1jV9KY5BDgLBq0JEt57jsWCQIIYGWpCRSCrO74mWE
SQyW2pxt0xx7dr0fwrBIV5ieY0fhBFoJN/WKIie7PkXVr5MNUlDfQr4q0MtEUSyW
xACkMEMmS1micQy7XBrORaszYd3yPxiTYjaLcEYkxDNDnMGsOatRyD3ojnbgAm5V
Lbehdl62dTaGS4RPzkqIyTf62vNewQ7AvBLCDSpCAKpzJkQaFtv81hld8Awgx5AT
JdSrqsmVH3Ylvg7z+KATBAPjCD/TFJKCuabknCorXx7G+oD3OTLYW5uFQlWvRTKb
9kUnCFxX59sw42lPuHqOaswF6VPR+R565ANCY4zPHhhhp+kzrDZDMBiFE2n084yb
f0aGdxOI3TJz5GI92uTlBJx18pwD+iJAw1XeDx3bZUu+yba6LqKW47eD0nmVCYBP
2eBm3b9fpM8osLz5o/vnohSvVeHu2gWJGie/yOC0UkV4sP4Hg+LMwimjpP/1js/h
hJhy9Pr9KuG3Ek1/Ptou6Hd0sck2qF4N31wdNIGFClykAFQyeIyiVhZckjBwOs5q
V7YBXY0sHH+lcxzb00JF/nzgqAByT2uH3O9T6i/pq0XttOWUMATmOcddeYBriegJ
4La2fUUXKxh9NRv3tVNMxZWBQoqeXCoZpnMbGmlt5VLpAIebhvh+XpXSQb6lS74q
k87vxMkPpj/56uPvnZB/Cxc2LyIyqmUC2uZpXqqfgrZw/lFl2yjTKAcEKtxNN+v3
3Co8cQ6Xs8uGfFFXkiZqLDvW+lAKfoaxPojl6aStxWsD7IUwrGgTRNlqEiyYa4nP
Rv22tYO5/H8vAc30Akdgj7ll9yjO0Kz+fRmyD02ThvBUpo56JnGOKZMXgynCvxJg
y6dRoQc708fWzR4qggykNw0sClcV9iidRTN95jTJjtzs8QMoCH7gFdDcesaWrL+v
L/f6erOG+xgpdewVC4T4fnufwMtTFwkM0zY3OV4LDXzc/y8PWvIouGY2P0MYVyXL
NC7Oun4+614aJTactc8P44wQCRdyWQKCr53ldaIkHDD3Tbq9co1UdQ4uuhzKxdlX
F6itzbgOdQzZVh38yqZEJHxB1hdE4ed8ESWjgQdnYAri6CPq7CepkYjl9uOqNv6o
I3HaUKeYcKuoAwSF8oLCSfM9fHnyAIl5BygLJpMJrI6IaEPxu9ObiLsSB+VE9fDy
kI5hIA9LgpK/BH+7dkdulciTbVEtjJ4GrkPytYRiUsG+TNpBDgLFZYJfLAyLQV6K
Kr+FFoSb+P6Awp0USh36MXeh23UR/s7i+lCQvHYX6yfS1WtY6Xop5hlZX/MOOI8K
JAZf3P4ECqY8hGTzkZSlurdFkzDLkGvLkNjz/YliHblTIEwCCiVGIWGEfk+4UrzP
dhQN4KIAZ66uK5bbzQTrq7WBDNkRsG6A2f0RQnnHbPw3SQgO9PJOW8SsEHfIAgLf
AzW0QT6U1CDvWyed6qS20stUWhkkqEziKFM2i0G77p4d9h9M2V9enyakD8noc7Dh
xgK3o8jp80me+5ll65yQRFpuHUa/nflqSCVrntxoN0vTMNCtLwA0sci/nJbaiO2S
65vNq96xO31VGcOJXCj27JGkRDhYxna6R2oCn4SUuuXh3KiVjQwPKmsoqhaK2985
3J9goUoow44G1jTEeKYtHz88Tumi4UqTfmS1QeVHuUKX0/mHVySNJN3rkkFGu7Jw
7Dpp7iuTUqaRypEhIbQb4LsCzLsQ0AVlpgEjCxjvDpDcLVA9BfNwNrXknSM0sd5e
s6UsEVIRTJnzgAZP1OxZgUqZAxCCjvTg/MZttvQOBhngMXUIDV14UQj7GjADtHmL
9RigWNQGrAzdsGsUurRrUVzWen9VEJTxW6hVKf1HdN0NgjRgvk0/hFKbVxdB2TJ5
dc+Z/PeXUrx5YUk+azUDOksPnQaB11Efr20gLUtsZ2F2VBIvexaw39F25LxjqIKv
bTRcwCVMX5WWew/KfiDax4TaLlUcX+802Cc6iqEFzE0PfapaExu+XeInbg4N1+Ar
iRMM8CiBTBpZ8DHRZUUcPj1Tv1Z9g02azA0ive3n/sPO1DWoMrl7SVHayTMo+9uP
KGSUaw7wvizRSHHIgm2n2npoBqf/fYqu6nKDgjftSIaJZaA+eZdogJA+kvkse5Lf
nbd+5CENH1kVcnJ4V7TV8DFNdA0Kewjq3dXXtPToKj6i/NJnpHP5TKT0A8PUfdaf
ePgVKGMOqKCfYgWq6krOoXbaFOjp7JqiVKmvKgP2OYoX19HDgOBgH71gzPQWakhA
o8mtRoW2gRUkAVwJZRRoSh++fXMlxr4Oj0djTU5QjiOS23RKDhuTLwI1RYExzYsW
3yHin18ZFxyiLf1HMrLoeT9D/d8ELFuQoz2rdPpxiVw6hCr0R7+FEOqtMTjC8fKH
UXb3TrvMSI6odoTWG+lk4ynv709jfY+iW6554LvDgXX9U74Cys/k9k00yqX8ZlPw
SZ78wOJ7S9wgbYye+nxn+T6Yf/AjpDe9eIwO4GB8EYhqEkTHH0B6jRoQZn0CDEUH
Ese3HdnsieKvDRtSWGJIO+S6W3lVM47TsIrp8XJB7maPqiLRaXDYzjQfL6QjR/ST
nb1EmUPpgrCis92J1f1l/Y5Wrf4+veE+Treoiu9jxqRWRIBhRtmbGmr0GtZe37ex
zr6OQNMnxVUaY3D7VuEZaDcnXlc/aOBItCmV/NL9RWHyhp8snbVbaHTavc+4MouX
0ukacq1EJ7dG0ZstojFcqC/n7AHZrB3NefOthOwebjQyDUadJ/Mxk7L6bO6h5kr6
vxWB6GZ8HBIoiWS6X4tzUOVK/vkNiY3qBLdkUST5YVpttcpt9k0OD7Y1jHuloKu8
ZldyTsNSX3J/RDgbvJuh+WNGQ9vzLadzCszfydOzPBOPKoQOy/k/Y3zr4/+PG4S/
IOZxNB7JUKu8SbpNvV8HWwf/GlwiTZezCDKgqKDMdyh71Mjfvu0DPX7BRXagu8fC
+kPH5fJdPoy50NGbXVIblLWgtQQcuub9jMHkO1w0VWf53hVYYCzum5NIbewN5HR5
AQXYy9U8IFaAmyNDYzAexPvBaIXpQZbE8tyJ6zcelQ6M3KEykz93ph5EwCpdRMQF
vE56OlXipkgRe6GuTPnGAQ+SfMF20eGxg+AQNwvon3dhUx1RKnrr7wZ5juFaUJrP
S72ybkvGMNM/gsZjWBb5aJ37BVNdWPZbPb3XZ3BMkc0PnPdSfczb3V17bhZAFoex
uJ5jEA18ESeHadCOu4G2FgLhOK1Yf3m885N1kL3bmAJgf0Wpbdh8diDHBCtmZA4e
wxlHM1fgtPdRbQR+jB/jIUK/oQsq/HpBtfK8TzpYgyb7tumPfEmHxRSTOUN09sCo
BhAgpfj65nn+lEwqAxE6cROirtAC7wxpeX7sSavzsudBHLV/7vRDgVMErxeoqJW6
EoGRZI8ZumRO1h9qsDBzm640VRJUjhLNpqwj133V+zFyUcTxHHKvjT3YDHkaTMrX
zEVwzbkWyLeg1eYrO8PhLmj+2ubCs8lhevn81rfTTEfxPeNncRbZFu9QP6dWnMh0
bAGBG/ItuzulurVCy4MUnfiNQtRVti9FYxYnUInQEyC54Etf7WO6NpChrlyHCq1A
CQUjn7qylLi5+2qBIGVQeD9AXxvx19cwjcfJStXM8osJcL+KOmBBboYmtm78Ascs
BBgLXO3qJj1NpuvPisZ8KaeNDi9Rb8a1eBzvDNwOxL8iCV7e59ngKh1vZ38x8i1v
68MP/MtO0d5TsAcqWe9spVBMYlpUQE6lbz4L5isaIzYFyXCPDmfwUxshx5C5taRi
QFfPQb0oLn+Tuq8gHBoq3gFt4f+hfzJ85aqHrSWwiPzogy2IlNVm8gl98EzUWlFE
VINMhhXoRBBVXUI8TTswpDr8Fc/pxCtcbV3M2xDvddpD3ZweWp2qlQpecpWuiG5o
z0HtgIckddQFqciCgvqLHOkHeFuf5G/OsxKmTfAfTUt/Bp+2jpJlOpQbl/JMXhnb
LUQZhyBAAmAW3Nw4vaPBnP8AipvTj5PC0RYcATTETLvIfz4WUt7YGjUKQ13xwhDR
DmX2ArtbphR333iJ7K+UJby9Kah0u2UWhbB7a4plU1RkgqzZnOQLFiZhfb1aicfd
YEzA0AtYjr9lFW2n7duooT5NnYbnpBWsc/NPSKWXmykRCaFEqwX0cr9eQACV4ZoC
kjxB4NxwU+/w4yAWt/3zY8czaXkNDU0sSHDOULaYnfHZViNIV/Hy0E6/VRJRi/cQ
loygKI6YrmwqLVRQfvFI9zbulPcXRnPwRusVZurhWL7Kxv4iPR4Nq0McTjdauXxK
B1lDIQ3NVtPZrcmeKAKogGyK18imDRbaL+bBF/Vp/uGpDB8IYA08xAU+04uRDotM
C7nRTWKDLQ6DdzVYuTqz1aneJln2Nd+3u31WGpt+A2KUROIldjmL200pXFQJFBSR
X3FEobN8xwucCCQrgDlEEZ3Fdzfd68hi5Aus6LijFvo8pXw6cJmY7iZsZFSjq1Hi
aIv1d95c73SDczuVA7mkJapvT5t6hgwRH2drQtxRxO7AJYumKmBfRy1OrfLxLgCi
ZSqUkWXFWV8zon0JHD1ocAfvF7w4To7pIYPugZOjCLpHpAq2O8L1MTLIiUrtIMB0
p6fw5N9YgFtt0mKsaBA/Vi+6VU96eHbvz6ogtePC0YsEou3wl74btAa8q+lDKiLp
ngKqn3wyD78Q3ef6zH7Qm1YGBIUdfLd2rdoMWKF6bggJkbqaHq98dDZN0hM9h9fG
/i/kCDOPGkHl/ZVBQfHiKP+g1IOP+5sjRKIFF5tLLq02+ZeUa65gqyrnnVb0Ut3W
TLDDQJ3RaMP6BCWEgpq/X181oDpUlZ470+Q8sQXS9rCKtbdiWype0fRj5ZPbQTw7
TuU5BJXUG4lGfq0DCB77qH3ia2s0VtjHDFQtyKCfjGhaGYP60YKOHvd8iSNWA8No
+03p5lZqc/N8NR2mDOzcnAC3zXoLKGzNvOg/mup7YMv6DVf53kdxJKfCX/fvUQMt
c74EMa0ygmn4Oi6Bo+b5ejtrs0SMg9ilzbxNw6QHP8/rFMYK2HzYhdBRoNF/NCtQ
JL+kQQoUW0l9sW0/5Cs+84y/0Y1+nbnZbrnV8sg15ZXlIxjtz9KQoOIXbmeRLs9I
Oo1JfaEOAEvYuAqjiDzr05djUQh1roMbkhooB2QzJz40Cta0We5LYXKDKFJj5FMS
J+haG9FRIFwy4wuuREQ6q13f2W0K0lZALiDpwxQCr0gUC1jviYJMJGvrifHqZt4G
EX8r8bqUDhMu02J4/z7xdofnoEQKVC4HMLJgsK5AawJTBcgHvu8CdOnRmRjUO7mG
wZaimxdZbEbZVSFUvGAAPEdhiLNNLcuLWRi9LGCzfp2KtoYWW5+LORvXEOzYd3DE
b4E0EF6oXUjH9tYafabkNjgH2tLAcCS6Tz8CIkJ5ACTRr4xONi4im7yJYtzSLhOc
04N+PUfD0uGZB+rcpMEwzYn9PZrOzA1q4ofH/x0covFGTCms9KQZN0pRvW2bovc2
WXrVDF5G2BSUjV2BG9baEnynnWvP2KLUWNd5XAyoeyUs6meF9BMw7tHF0nxkp9Mo
UXI4bwWsd+cXLS4YTx5WSv5vpXa2mStNh4lbyz+zw94L1cHDs/OkxentbcG1mfI6
37YuUUVCeHVpkl13XKXbTyiMsxGOQRmBhkFDsw2MD3OCn6UUNgOWZnBCqNd7xRoh
HpI4GCwNnWIVp4G5NQ3JzBbxdHIh+Y5Y+OOvlXSZH0oxDLYV7KdybZ0oR3kKXBkT
ZcbYu7DHi3MbI390ElSdzm6DbspoGEuDyMGGOWnZq7mpVDA+xgJcJD6ePwQ5ZC72
/7r42vXZBCNcxzq+fmhOXHsJX0d/Ypm31tlJOmp97GPAbwZO7cHohbqNrmeXCapz
93muyVcs4Q96eCMZJH1DlJeU9ivbe0EpEmjOwWAAWwSsz8Ke02FfgfY5NBgt1QvO
xHrrFCN7VGA39MNMJ+z/NAtLleQCq+sfrrwGsycLGyO4CMwFBX3T82OuG0m/Zt7h
BN0dfjz+qyWwHHuPPEyZNnaKguixyg5XhAsEJBRu73AO/9WoPQXkXGHs7yVbqXok
Fce0hQ/whx9S99kJEKY1jH1ObOaPjUSWWE48EJiESf+VZQgU/9MqNEjw/gP+JPB1
7g8pUXakjjrCSWvxQNwzgiBJ2hBDchRHQ7xhXdm2XCf//IS3X+wfo+jwQW8YUlyA
C5XeIn83DKIXqMZ8cWLgBjCw/qtRte6ZflZT5PkQsagtkBf0HW6XUbpugvkz399a
rcQhxDPM/pdcewfjHy4rXUA7mqOHS1OemL6Sm2y5RLKkelQxBcJc+KaEmXTSc7ZZ
OcYyRwZuQUUtrUsbyHATkSwX6i2SPP6knaNoQneztd0muFKnl0l3pRaoDX+0nK1D
TOUF7sz2Zw4CYoNrV/GMjxRsag581Bm/Qi/Y1J2EuBQOxY9OskwriXbMQv8FBb9j
r6/hXj3tVWES+Nknrw960Xi9dwL4uYinPWYh+bxuLp5ot5BRrK/VCYHUz4SCRojb
uN5/VfQU8lK5cIi/mwFXzyFgUfdTG0SXL9cFyW4cjRflm6+tFCwIwNYSkYMUUwph
7CJNfdP2F7igSKpODEG/u+JSBJ5H4LqwqPH3eOMXjbNFx4rDTF7yri4OEBqXYo03
oL4Itzh27J3B9ALV9fcWaoIhgAqi5zRWWw4wv9NTWy5pJNg9YzpjHU+h+s0a/+ix
60Vz9xVxpcaosUzqsGwEcFnJyohSMjYs59HI9UnvNl3R7cmvJ2u7ejTh6/Xe+W3C
gCarSbwSH11uaq1+DeCFrmxdLu0VB7gpertFpAQS9oimnnDiVINwrmq7jyz9JClA
QSBN+eZ7qnuGz9Aee2KLFrcrTHMWTjbJIflKMdlGdNGNkEHHJHgYTy6DGt5tw4xA
p9SCyrajI6Ax49UBYIkbilDm6/Ok3z7mJWtpw+kNKcbv9+d9iU+yIrwPyDeUhgSJ
kewMm4H4qYHE0+d8IFRiTDSg2GfB8AftbdUtDWQ28FehA5EARDwf2wYsn4GjB2Di
dQ2b3q+HUNSno0ol8bTfCRXXMxiWhiATsdeiNOVt2FLhwK4bbwUBpS7med/yIywJ
+BNF2Y/DWv+rixboISfYSwEJlr7e8D7AZeV4rULhIAdgWZBupZvCPquYMI+N0Ss4
fSTM6JyAhwj+VvB7dgfVs5S9sM1C/dtIwxoiV3tPcjtGe3vZFjiUlG6DFp6jL7/1
s9Mwd1hLf41ONOkE3A6QW8N1+nAy7PxqRYOmQyu3n6l/dqvOXXLCGbBUeol6SrBX
QOMIbPAPafdohz2XlyusEAS5wsHHHz/PHKFs1tpygpM4OZzDgl6BM+NI3v8TU6/z
Jb1b4+tmEGwdQQ6FhPMbQgQ9wueSYSkr5/hmK74pxkNOV32X1jFO3nKxW4pM0L9U
cwO5l76Yi0XTQFysf1C7MPGNfNQpYrW3+gP7Xsbf8kpyvsEQM2UGdpo06m4cY5yL
Id2PbfyekbOcJZoHo2GOCUZEsj0J5Z5gFi7lF3yyFLLjDwUd5C8ZOsMqvU1Guxyo
LpsI4ZMryjrS0r194ojaooHCKsZmq3Bb35oWPszeF6t1yZ5XmRUH0eg+JtbgT+fM
oPHyWtlBL+NVHnpXU384KROmGaKsWQ3rI3xAjeNqoameI/8VvcqSvTi2xANG8+Px
E/9VgueSZ8M3EOQK41GOmOGwKHumXqxytDv+0x5ectd3kFIaRNb1vRxLWjTpfxsI
zzbGh6qtXSubfAVpVvFNDRKYDzcW5SE8jpKQH0p211d6WQ4Q2rhAV2ORqjB9jP2c
y8LrWAf8u5Ypcxfnuxz0polBYliM1PsYzQ0J/cjbPIayUJGSaXGRQdLwz6ZnGFGq
VFZKEsCZ3aQcBIJhnAe9kl3TbcNan8zHjVWYSxt3M5zWxDhcKHVeJz3le7sDS+Mm
RWH4Y6CAlQ7dOecgnqnBgFlGPG9gYj8O3DM4HGgSYMAIzryUDfvvSka7T8v1F02x
yvDmXYi1QIyJwBj/pdyyAzDnPaXVhfVmt0gQh6tChnV6054L9zqGmIVwTfJ0hSB9
NLs4XkVwTfaYOqZA9BQz9S9glWlTkSAHXLfLToIkUnghl7mJMAs5m3gXEwyMkxoy
JYZZayqvOEkWRzHgkNPvO0fKApS3SgMRATnQGX1nDWrAbTtWZ2y4BtQNO5IywJyb
WLk4Pgpy1bu3hMcoVCBBrC3ylWOuJV2JRs53opmIXUXoMi1lTNrLM7XHyl+9pu0L
oI9yfZAHk4gq2c1nvWe2Vobex+mk169TiJDifV7TEl1Dm6CzrhQKbtvf3Jl5rDPa
XBfRbCd4n0uByTr2/vGMXOJTDWAPMxBxWOhc1IgzzS00bcSl+XrDC+ISeaMbNhGg
3vnRGZpoQxMTmy2xeWoeFvO2jN9XtB3t24+EBBW8hZKfMuw41cqyerRekqcWrLwd
Nix/LL6EHi+Vnf0Du/60i8kLP2S43Kl+LGivLaGJwg0oTbflaG/EdG7qVAoggMxt
V1b/ccUwnnWSBAXoVgnUAXi+Anm++caCdvIrOxlf9i36QT8cRFWawFEiNNr5pjhE
IKBeyf7HJMTdF/R/POntVj2N6U2/Z4+ip9QlJMVM3RXHWv9V5gSsERN/ZIyFUnfn
rSauFuliY9CyL8IOHNrlBnE1qHS1wX/LozxVqR1pAa/tqGxCFSPc3gk5uAFOHzOq
KIoz1lbnuasHkFlxAZY9ZhltbnEoXXhM63AnXnDSvWH58z6k/FvafezPqP8E49Ys
wisBz9BqLL8eIVkfAqUzwTKCS7BATfjQ/SGKiigqxuJ75j+rBgt1H24WdAMjJ2yU
nQBjY4g7xGEWKG3Pz35voHk0EGqJwrkE/sHz7neAlHOT5v2jRUgEJ7iQK90w8mDH
MvY9zk1ajtmYxb8nAW7tZ+nbnb28UANj41oK1lgaSUkNBfnOSUTEEGJv8LppBWpN
XiywQMXYPUOA6DDXlnBheTtzzVPdPz9Sbj9y3sc2i/88HKHAJUpL8y8X//0SLYfd
CdvnVcf3f7KQWB1WcKbViYw33Ux1+eIuB4SoiQXuOHFIsgdyPxEx7GbpjIznvvN7
TzU7av+jMwNRQ039T26/ZJUw10Ysxd200qeSP4TAzCT3RWMauTACM829SuDSgsP+
OgW/XV2v6qxQmcWvrZS/QDSfyPd+/WhVRhO8vwCquA9dFzkKfnWFzMGci2R7YCO4
dUQGiBtUa4qUn1t8W1SlFSFig1VHmijOufzi35sa141oDM16gsFpbACeziieTHmc
GMmeOtIwQs0qWHv8ung72kxeNetqUQtoOzxSMPsWVoAbDp2Y1MbIu4UkbHJ2XpFf
4le7lXbfvS5kz2lCTvl1PwtBF1Xp1TnaslITadEzTEK/04U/e6zpIPjYOBI0QdsF
Qqbzqp1W8InwqaC1pCDIbyDWYnyGhb3+ZXOggBykABTVmkoxppjLBIHtzMwtYZS2
Ru07vx+TiBMkO28E6MnWPQNnQZZEV+nByDaoHaN8iDEfzVfj/LgFV1Yx/M7EM3O0
1aapDMk3mGkXvPD5FC0Bu4MCemU+YquyOQU5V5rrTN8gnigFZGsjIemX0P1WqKsc
cnPMOd0z6t4TFAWUn1UhLuCFkWm6EF59acyn8thLcm+tBZvtbbLX1+9sxbIRFZQP
pXXzS/T8jEKGv7zEzZlp096zH0O7LVsdrPZp7sEvkLvJ1iVA1cjD5/j7xijlm5jm
eP6QiYyotWcsc7h9xicgvtlY+9csZB0B0H9wUnbikLvH5X7f5YCPVUfH9FZCNALP
mxIeSa/cOHTcDVigE1tZco8pEK9gmJ9N+mBXluXu4AK7jBNNSXzHGGBJ8znsl2sY
DR3zZjJgGqYP253gzTp6QMEODdboU53O9KBtj4fOdHqFly3sEFXsO58ErjX5HVHX
eOnnNbneX0rx1vvqRFag67OHKbHq6vNi8vwLLjWtHnz7jOhL9wrpFklv8ciiBV0e
KdUT95TuAQEPFyB/imQ7c0s0Kvuyxx8NLfVX0auECerVP7pbG8j0qQDTTaHEXZra
6fLlQ5rD5qB+dd0I1nSjE2naIBepkyJwsYu5hWSCDMCLmyjSAF6ZG7ZYYbPgIo+L
znxgCNFgTSnaVIUc59L2HixGsNej+c3rsXDMvISNT5df+7882NA1QYkDK4IAjoA8
AmShugKbin2T7r6uD1Y3UnXJHUVUcPwMkAPsAWtcMUpsDoeVys86DSub7qwOg9M/
eckMShfK2mnKeln1z4RwnGiHglK/52/pdw3Y1DFieH21UPaV9v6PO9kFennGCN5+
v2j4hV+MFDjCAlqgCwJS+OIiY8ShHJEHqhz6okc/5DKtk4VS1U/W+yZLiQxZhDOR
nDwlM5BNZ+6idCoEo6aebeWd2RlFSfRIEenML7dERcWHJ15llElHS3Z0vDzAPyJH
bKrkdXF/yxhJgZLZi2OoInx5dAunO37Gq+FfUopTnVrOR0i72hb5bddJPQYSAgAh
aKJNZHgxh7Xsujiq6cekNgq3ER8aREBSx8PDlOt6O01wf3lt2FOMQDGx8766lmAG
z+ZutXqY49l3GHkDNWRI8xoQCinwlsNxeblawRrelrbdSdbkV99D8GShEgJCh6X5
nj6pnpP9z8imHSL2WFv81YJQCuCkL3p7qWxSZdkGeMzbK0UtWBOkdLzXwm98IM9P
T9Rvjajwz0TeiTzcyTZW+29EPBl/gnXb9HIKXyqhveag8tL2Gdc+XPijM0YwXFqm
qZoo0CPBg+RsMryCYO9iQvPwa9SSyRilxyBH8dgHov4gE+FPdk2JcAUXvvGTvSU+
WlLzMR9vVlmUh1rzevlH26Vki4u1r7vnoe6zJGAXwO+XRqRgP+PYxNTRfR0vXk3C
ckquVlt2/g6LJOdBFGviTd0LmFRBOIsMoQN9LZP7IR37TlP40ynjOJhXwLNQrc64
fa2HQHFhMHyUjNqZ9XGhVOD2QGe/zblED7SkgiiTnnB0IUX+P5mucYO1O2yWTi6+
D30PxSfcGlkCAB2Lr5oxzrh96zqu3P4Lgm7SgDDLeL4mP7smbC9pClmcp1FvQ7uj
5Rha4YJc/xddN8Z/BYfWkhi0P0m/i+WMP2S4Xc8lFDPbG5fHl9/hHDsmzzR6JQNM
7UFar6R7BgYSLZSmkl2R48YUD0h90bv3bNPQn5Zc/2SECfPRfJ7fnhvSgFMhOYwm
ZJyoQM0l1VRdLGYMBE8VSMzF6R/Ksv0t4qzft1WlDy2Vo4DadaXyLcQ1S0eFQTpC
aBXdeINoMXTTj9upZb22b5HupR2MbCg4o570plZoHa5c//ba1B+QZsKxejlMLNAB
v47qXgLsCPfaYvlSbp3vLLyo7Et7dbfKDXCobe63KIFdoF6SllrZk+pFmTf8hYHQ
HdrIFgrIaWCb4f+9Cm6Foa+DPrf1cazRE+vmzmBB481QkDJM59nB+dYI7N/Eccpg
YpbhjJoUKCOBid9HZwxsFY5XgNE6bdnKVqBrSOueHWocf/LkhnjMF491Rf4lVAFR
mn/4+ch6X5rEvC1p+F8OCTFlnKkoGrzeAKjt8iiX9o05D9L01u0dBWrWfZr0UuZJ
iHwkr9fZGcTaxxQ1dIeQweDZF0RSxHkYdGi3bM1kgfLOD27FP+Z2j7qmax/x3vnj
QFNjdENNDCEQuEjfsWrAJdfid+SFaFnxQIdU2TgQRF2pmWLhiVDgTJmV1AXRW8Hb
//GXw8iFCoEjB9IKmkfba+ChtMGNlUzrgTeG2JlqzenJX/fwg6JCUEHTvyOFXqZp
BdF0sBOk32h0n148MkkKKqCnCvLCvHHIcHFynBLh0pC5Zwp5x57qQCXMsKoy0xYl
ZF1KMLcwfwUrreuE/1Nj5rQfkr1h6czNC9r9y6rj4HEEk8rfYtyTEKc2l81OH3po
q8XC3TAExQeJE6h+JhIeeB+US8wR7S3Og57Yzg//JQeBR9TS94WQqW1cVZGCcuXG
rApuj+58zryLA84XLA/UMB6AhB1KPjYh/4i5vwtheBbtlS2D1iI05Ve75Is4NwB9
Lv/C8YVoqfqCBPaYUMPQ9/KuJXkKRvH4+hBdDoTpP7lCHxCOKvt8qp3LWXEKvfzD
VOlkpx/rcAlhbmzZG0rAU7RjVSnLsBVj8s90grgIgNz66hYkR/ZdBlMZi1WOp3ad
kQdVzo2qUk8+Jd6QoO77OQuXuUbdtcUnpBfM+Jod5yZIrIcrRi5/5y6+pZk1BxgE
NPUT+K6hBAZG/zY/Qxheg9bjb6MXOpcI9Zd6FFmH4yhjN/jgfUkFTKrHSY0pSOjp
SlemCaWTp0x3R3mDPUFwE7grk0uubHm4zQWCGED1c8it7Rx11dry6jsC18EDpzDj
4rx6eZKmNSVU5Ban3P9ioyrOhuQ4EYZ6Svs0mx6FoA0A1pCbvu0Ercr19K7T0EiV
lI3XnrRnLohbE/DdW/bZ7oJh1wZoq9Mu5q5ZEYu7/19XCmkkoDYd7iUjgOmDLWMY
W4358y4Eq+4xjAZvSPedAno17FHzdAymYeSzerrtNdXHrmSOMw1X9YtI18Bxeok/
bM0wxrc2sgda0PeF4CyZss9vBYgSaKe02FSFLJ/SR1daG5zfrsTtXoCY5FhyZGWW
4VGc74fLsI7TNXu2dFmxpDi0i8gToy8RPb/c+46KoKKV6jVODvkmPkY116+wIxWW
C6hbpO4EZgdEGbk64g17nh0TFwUdf3J4GYwu2G6GbJPwGnFX+3MqTT0bQH/dPXYu
vgf1c7KnopbOzwT1nQIe7D26h0r1GiUbv8qFPs0TcEnKIVs2vn4RK2xXFqTYQrq7
I5iMZTNGbKOBQ6EpOUbfbAxOt6t24qhhW3vfeqc6QPVetxsIMliKI3ApkQ2CIUoz
eWdsA4rAKYbowv+DH9uLZhQriviQHr3PnNPVSP8Po/OCkez4cUhY6DUh4M5VlMtO
ZVCsy7PHzQ5tJ5HAnYCLsD501fPIKWVm4Bd8GsbWY1vhqAyPP3R7rZS21pL3QLn1
HV+EqWyx6vfDsH7aQ+rdN6UEUOJ8F80IlLMbhvpJ8jOlmfb0TL7r6CgE1nKwtTP/
8VX6A9zT1DnN9SQ9l0avIpRt6fEKg4XQAMrqFYIn9U75y+CxfAvYL9iPyXxKJZYc
ws0A5xleBgIMGEy3rENROT6FrQuodXlG+jBRSL7DdjC5Na98EdHcaEWtJAqA6LfJ
wzLLBQB5S3BMOvtoGQ2lVqnF6N35w+KJZsB9wo+Pn/mQF9I3xjSlzvWOIJkDLqE5
dgClrZFEzZfyO4EDkLUPR++zdFMgG3AWhOKdTDos/VNPrBd13SE8efBcQLOhVEyM
OeMjSnO7PPqwXqC37xmp/QOYmhyvx6ufS247PGNhsrgCnNFdY4m8YABkuv37bx+h
4YP3bLMPsP/VChHYEvl+TJqdALlaXyrETS0TTK2GhVHggFh+vooOH+d5gRvecJuZ
iKUpbAhVqHXSsgH7x5oWyvE/aG7zL0boVP5iBZbx3lVgYZwwOvFbnWQiaSqExD38
7J+ubjatX1o4tc8353RuM+pvNp+aLmtAGaqCl3El/X3xJkjfobP0kFnCmahn7UoY
Is5HUvam80B6R6Rv+XklK6W63AID78L/RmrEL6Ou6tIGg184iODJdkL39nH8BfNU
cc1IW1L+S4sEsBRWSaP6tzX2/9BQiq6WjtfH9tGBWp26zz35a2OFgpwkZ7OVxjk1
sWwQO1l6Sf6HtjFgeLWpi69nxn3TjqA/pivhDYUupWllowPO2rTYYmPmfgFP4WpP
go1eq0CA2c/BhDqIL5WYDc4lZnHNdaaTlpiBRwX7YI2ZIfPIP2wW2rm9TkQQ1uZd
vWJ6K75E9PTsnggrMhUNwW4Q6joE4nqeOMHouztX5V1GnyaX1QXtP6r8t2dtS/jW
XZkJdg8phuxZcosYxumvCCJ1noYaH7aC6vax+vMKqR3RSOawBSKoykU/fcez2oRK
aPwLO/TpFEKTSi3Tw4kfkavCzVjBd16ioyzVai4fgt5Q/Jth4hP7rhxXhvnn/E97
az9iGg8kilywRuos52JjDeWQ+EzSHghweqxurA3nLRTN69r+PliNmULmHj6DchWt
VYUBSTmZuuO0YNm+i55R1/VHlm4xPuJBBjCLsqsowJWZJEm4NdBSOgZfbZdZO0T4
SaZ1+9CB2jStbtOFZyHwP4dzCyWhmm8CrePUi2kCUPeGMxpn/XCxD2GnMQX9377m
dEZ2TtKVEPjdxTsicgyBVU0EdUVMb0leVv/f10361oeYdT83qcNaQ7n8Vf+SC2Ro
1wruc67BmxLvJQnBd9NjofvB7aF68+zCevBeboh51nB2b0dpX0IurzZdOmsz89UU
+Cne9jz/GvufYyUOn2/WF4Y2xaxrc5X1lAk6BpNHYA0UlSDATghac/07RgyEQ14S
TfvAoWWdWZpAjLO+YTeea9zD55+i/tZIgvsJnY8mK3MV0d4xdj/5fDPCW1CXULy1
Q1ScCLXJiJRtFpMa1GWdv8cOz2WmeDDhKya02+g1MoZmtHySlp0izr7WUl7DYKEh
/tA6NmcHVb961zuSg7St/phYr4vJzcQGhWCfLk9JAFhLnQ36sohSK+/jYLslwdNy
Pi1StbZPMQFJGXtgVGmrOYKeLsSxBh9RRRK2ZZqCWZjzxOahh/TcZ1L7bCslsBUP
CMzgUfSC0kra/XIE149j59tIgUeK9W5B8kFJ5c2EYX70dkjF7ESYihEYN2/35j4p
7ZCXLtnARg5x/wAuj5daVuyyYrrx+C64FABm1QIwYT/IwutV5ve+pij4BR8CAeQz
+y/enWIchA32zFKFPhRL31YrI6JLkmNHRCAOsq/pWP3Eo/cDbMmeOPY2gzDK8DuK
YUPqcWrvN11u78WKsa0bUVqYpJibhKbMIr6JKb0cAR/rlMtmJNFldZBEcEBf1nap
RLJVL2Q4LEeahDSsVmHzJVVrwjUuTZPZ6UdTnfj2DfJhVDHlyea2eu/z6VqFTH+y
z5olKgmPUyP9uR225SMk7YDLlAYOJkTFDqaN/D5mxqT+n1g+TH05n6+K0ukYxORC
tBwZO3yiUn4BpUQO1OEjbtTTEyQjEtGyw6Qv+2pVv1pELT/qtGVXMrzDrIqeXlff
8v0Fcl2SmhNNYeHvxxQVUWk+O9QtaAjHlpGO05g4HuGjKP3o3/NCDAFvidZvJQhc
mALktbeu/F4lgkx0Kyzq8o5u8qJfoc2gvyodWD8XRYzo/60oLlx6FyAPqfQnyO9B
/Z5psr7VJC8TyiTvzmES9XjM1jh/qymlBAWQv+EcQsHmeUOZfneDBwvkMFJ5+b2K
d5j0tx/Th/Y+9Zf9MjPFd4AZLjRjoUbMArDsAYnWj+bB7382gXOHjGOPvN/VBWyF
OY+kTU/9iW2H4jeYPxRlIw/eQixXLi9E46U8seJxrLkKTQn2iO2pd+4rqKV1SY4u
79jYZ7tgGJZL+obHpojjfva75BccldZQOTPyU3MZWrB4PUD6+6XFy6QZKzHQuuZV
zwMmXmoJewTYffBLU6AWdSjtNsKLIBmcKSf7/fG2C4LUsCoLN3VUsaR6KOm5Bs/K
IbqmuoBnj1bTpw9CkU+PZ8pGXnVowmMJWkHrm5HHXMoh4zAXXjSJ8lAEml/sx2Fp
R7zvVnsHbIPZZpVH4H0bYcgJ+OR3k4ZfQxMYz5sWAhCDxDhApD6Dn3drp0jFcfJZ
4AxXyVRDB8ifiEekHIDPPwlwoyzH5d/O23eBdeslxZF/zuzIt5987aGXzsgOCnw6
A+o+pMzj62q9/qUgkeRrqjG5PSCAARFmLrYTFItVsZMutMNLDujTeQbnloUJizj4
J/cKvT3LwLN+D/qkfqwAnifYeMu88e3pCiX++VzkC5bDt2SY2qTg7xm8b7HE71+E
KfkSHS45cq7hhUthiLExmetIPAEIAKk4/1W5TYnmsVfcjUcI9aM1kQOfzU+oyGkP
UjZEUe48CuvcTX3Z9jq6nftfdTC93joX9yYd1HNPJA6Pn4ZMuTCHJ70v7RvxJvfY
lwHZxfmpWrLL2EAnV8se//frdxllBqjVongGmBLIgM51ZzXr3SjTsW/LRH7V+O4a
mEkz2K4hhwer7tQeKdOq6wVStO1ETwVfdeMnu/Z81Q8at3Mdm4S+se3l2GQJa6G8
utWHQf2qm1MIUd/i2JeLwP/bo8eHV8jlmeQ1pTTKfrF/um0JrQX052rBodx6Re2h
xw0SQdf+1zj37babn4QXTTW5yyzdrwRbRuj5M2g0T4vkwBSGV9njTx1QlXLq5n9m
tGCINHmLd5KdCgCva4GvZRqYLbZGJSUefLnz4GIvkZR+xcwTPmUduzZI9feQ+2rK
gQTEq/1ltQ2dtAdke7GRyGzfGPMbxJbt11LiKH2IiN34BPnQQ+ZgxsOp92eqprKp
yWUipFifACVicq5JexkRwUz2RlhIK5LGfU4j29vKCAYF/5SAeZY1IV+UL/zuMpN2
iQ3FnPSiE03E7hRVuznzcXHVk8LDxjYpqJWgr92Eo9gkqj6/Mp32mZMUUykDb8wA
N5FNJJaDxuV2W77QaxUVhwp1HPXmtm5/lSDjwsNwWmA8o2qeUpgZCsMbBainMcMm
0lQsEWO761zyUu5sHFelJ/DFcY/xGtsRfgqtfg0OvJZWJ3xnWDtqzuIdtvt9MDgj
JALsYYMuVflAHr/Jghud7KYeqae+RH7X/33Jvo02Id1g0KpERYicYt5gpE7kvsn1
WIcLWTM57l2BW/kQBetswPTqkCo59qPSwpMPkLZzxomd1XmbfOZWAfCTB0F5gjD+
glkL4+R0WaE2dX/rwR8On7tVUJR/3dPvC2JyKZF3hqxcX8cNnk/gZn4k8UJRrMa+
gVZk5SE6883aJ7vyAfGZe8jqzhwoOo2b8ZpuihHcLgYBlcyLSGqFCIigYZLkOoYc
VEWjLoN+F1F8c4BuT7Rwj47ZUeJLW9m7kef0Ur0VCZ0O7/b60oFfc+H+A8+SP0gx
q0cWYE+GVHj7naRzFk89WoLx/GxbmexfSmZZ/f3zOewNhzSXv91U5NA3eXz8H69r
3AFWs7tz37GSaF86nX2p+G3aon5PQzZCZgPqM8IfmMukgjRZ8df2m8qPDh+uMvEn
ylzo/kNCeLO5Pc9egV1wP4/51YSdhXzVwS3FVDDdYerkeWZcEUwR1oO4x1ZShhN6
ZknodSxwEKc50nwnJ6+JC9rOQYMUe1V0Yw/H65HZkRUTiD5BEP+jw9zXjZSIJRkh
PNKsSqQ6eCexq4xfNlK4y+8QT7jvD6SzOIXPjDbAPpkbbZeiJTI2Zu++FlD9aBKz
9VmW7Sg8GV3vu9IBQSbL+9FedukKNpvJsvjSVQK0VsFCLDzGQUJk8L74GTqYuLzK
vYaxQSJhQ1jQfYZAI2awelflZ45RSSG4UbveFbSv8ugOjQ6N/77JSH6mPKTQNefl
MmYErIkD1LJvlDbI51OTQ9F4GP/GyusUasazcqh0Vrt6P2Y0WadRZdVbsvp0nYKs
aXI/6i5Z4D//I1uNWb+iCwUvh/LstZELjtNM8UTnp1OzP96jBpbRXtq/RZzLI+9M
YJ1WctyKstnqhGQY0hNrfypoXF8AbuxIlhRBthBRAHb2B3yM1KauItsaDKVbtdpk
oqV1G8Ltd71s8K6Rhc1o5XIfJWTuzmpmeDo3nNxm1IpGIlMcngTXv6uV43zcKf6L
+x+7XszWLmzOetUAGOeX3lc/Bt93G5hPxh2b4hMqmo+C8C0Y4DdWpBHTA+DuGj7t
TnqsDGqa4mZkbEvlHvw0vpNKOUyGuwMW8vSsUfUu2xu1uk1eG/TbiE9sANIgxzG6
VQw/AuKdP6/Isv19Z/oN8HOl+3F3fV/YAyS631w0VyXcAdzNHF8PZVtcmOS6/WY3
KgCWGCtB1sbjRxOljsM1R6XooT6rr0Trwmtyyk3M0QTVUI9o+GwFIdh1KPkZGA4Q
CgF6Z7iOyCKG5YV/8EwrFu6UtovdE3lpi9h/GAIoo92RFOMrHcUNFM5ef9hbQ1Kj
/+/eWOjBfk9mhG+QBOmj8b96WfFlvzNS+NeBX3HomCpTBD7P2kunndk5IYImV3RJ
39vBxTPf6AqaguZ5Z6Z10RyxnCpZX2wCfVVBXTCWcrN3HQ20r8tcMKXggqYr1KkI
FSVADDywlBhWyrqJTfQv2hiLeQOvVZZdd6Cro8uaDKQxr7/ZrF0zxRIe74qpyZeI
PiUisRuobqPe+DCt3Go8DAWv2kFStMoAPWC+7W8ZdQMM5sf5qlN0g8sf/ZFx5Sq8
ZwZQ6YeZiiCUUR6nWB9qLfp8yi/UupGJtYOrxB9A6R9w0FTZbhtKN4AENgSVPquu
OPjmIi0BUBY+G+0kRvL+bxWbUCHowc68SgjL2gKghDxCaWpV98TL9+rmNahc877G
zzHucHx4xq/XkhWBBRfbkTwhoPpvxiabXi0RFB6+1A8T6gFt9jO5hZYx+dnOPvlA
s5SAVmN5niDDnRgVfoebYP9aa1Ta5sbN1J7FkiOakc6qUbGojQ6xBa+HtLwx3DWQ
50Hbg+iMs1Y6dOh0Ax5F2i08Oao/SxuTw5hqnATqnLmgWGBZBvK4Wl0y+XkO5QFu
67rMff6NnTxBsayichdDXbE19n/g8KxjOWNwZBRojE+p1ncQz3yrRf/S4ni68Tqv
mlgOmnS6n8AlCC5OewRuWDYRauH96PICVIT1UctnSvxVUdc2SZShTS9EWdfOtaXx
aJUCzGaTeE0Q00llUy4Ea/WFEAVnFceIq4Q7FmjMWHxgqtZ2yrdeE+luk3Tqv/A4
ek2SSaU+kd/kQ3ZglkKo/2Mm4NfAyhvs9og23K2bH1rns4lvFfixQIQR14g2G0Wb
EkCM6oWMaWnXu0mAGUImGaDYXrH9GljW8HqtBlfve2RuXcDfPmyvqM53a1FhaVy5
ICzyr6N9pHI6Z8mAx4/H5DmPosEzggIdkywp0sWb3v02g57Gb+UaiavBrLNfi6oK
hT83ZZSinUwOEeq89f3UAVC9P8ovJ2LPgiSwd4+cKTNUOzMz7g4AD9vTubTRpcJq
8CaX8VnzkcEdt2mKHEZfDFo3HaV6BbczEDzVF0QjhAznjiIPDqz07zzExxLvgKRH
BbwS/T9rAoF/cEL6SyJwH9Pla+oVM3c76r7R/viDA1J1zWSFsrjYBmAA2JUemmWK
Qz07RYWVQbfe/q17pap/owoisFcdLs1VcqBWunodPek+1dCRnmo7OvhebeKKtqHC
QkCGUOi1GTzaza1S4Q3SrcIGZOdsCvtfrU1+9u31OFWl/uUYoBWFdNm5GNn4xnBk
n3/kYpMj72YN+KU00IcZWUkc5geRreHofqXQ3xGw6Rvo3oDNeHbxy63Tsa7Fth0X
qa8LyRzKoWnN/XX3T6c3+g7eXv6LlBY6rVkECHlFlAVodaPaCR1uiPAkZbKHrwte
/Jgiz7Bi2zri8gCVIh5vkcWA3UCbOcsS5F+4e05ql6lN6nZNoG8q71JviBgH3W/L
w1TkQ7AuzQD1Ag2QDDaa0aUCXsrGv9ABWo+WZHYOZvbEQAVz57Cq61f0n8bKIIxu
VGVSrXnZt5HzcJAa49ErhwjQteZnMdR+osjnxYbONksxG+jZjjcjINTQ9BBCqSs0
RVcKxGdiPP2q2nnYRkrBjlDc39xQbahSXMm5/uTsKdSkThpjf4INVZYmGU1TPuYX
NuFGNRVwj+9gk4PZ8RjyUiNvvxlmpn0llE4lUE11uucabogyqeQkjGluF1mQmHq8
75jJld+I5v/9dtsE7Z4Xw/56GylMgLDi0VYJoDQHfCi9zgQeBPnungPONVlpeTM6
O3xSWvKYsNao6iTaHfqqhPUhJExyKFOEzwMq7k2F4ad0PUfdFowE3iX/B8nf/R2I
SXaDERtIrA2A96vY/2KPlfl/q57d3wbwI4S0gBsVwhN/nqzdWazfgatQvzaOZTyW
9PrkLf0gau1ix0rrojQrB0WzygtktvQukrsY6+NqHQMolZyznH2dNUXPcWUc9lMs
OyT01IvUlFc97wiMUDaWLaXib5ijtQMzwEGBaa7tmUKx1haXCvddGD9KmbvESrQ4
vAaryREyr22i8ZI4FCxh9Za2BM6U/ixT0IAbtuGB2LD/TaYSpiHHJrfDeF8nW876
2lr1hmeLC9kAjY6sjnOYqdjlYV8Gb4KEqlDLDNmheudO84/flmjkDkt9h8T+QqtO
6zedH42bOs/7BNOZDLOUZk0dvxiLXKIiOGrZeMrTPqZqlRwbjb9MAymuLaEbrJaV
7q64GH2BMex0TlknhMw+2Xtv2uXwGPxGmt58b4Q48g/ANIkg2im7p0TXnpunQN+R
1SCZERw9v5cXvBgCD0yGWplk7ldeceiZeTrVhGpZuZe7iqG2y1bOsyX0Xsm5wCuJ
+rGmLZoHxBxoGORfVRPaM+q+I0jn7rH9UvRJakbzBHjlr85VRjWqMT3KOOda8n7+
Dr6nv4UtOZTrQVTiWtTfxCbidq/EuLFWr+EdAH+04PHuz9EJ2USzNudsDqiazkfZ
B+OBieAhP/kRZgvV1mmc7XlSBYCZu2vwhBJR025+goUwB+lRb2NnGfWJq3f1qFq4
wjTHtZKf68OlXVlZHzGVL8UYxBEz5mK1PvdZofS4ae27fU6BoX7ef5oI77fcaRvf
Q5nHK3BhB41fKIVR5PKVeCbLx384GsAeC3jWpDIz/VrciC41YDCXTikOcscXN4Hd
eoawhr6OJJPQUq6UHHiKGkLjUvK+dTxZ16b0fyDRjm5YDICrjTPn8IVSZYLuBpK4
ZafZDlUG2bAWdtDtt5az3LFmiAv2xgwY0aFQMNr9UVpSyERQLeJyxLKV+Bmbckq5
1yjK3CzCVPnfhoDIR1xgr3q7QuCefkQB/ZPTKULcZJ+Ue2L52ibIOi5b2d1lu4C+
CLhiBJVXWMlxhX9UTEwpCm+JvNvlbR/rPrsOoH1DSO8ADBQTM7qGbm3TKaSInshp
rNMBYjCIJ8f1WuymnPpQm6gYft8zSrLPOqUzqe1BmHMZUQSVskYDWTyYzqq3YS0H
Jdm/a0OYXGmpcGDpH/4TTEwP29KaqWsfhF0cevn6cvEGyKbw7VnmRqOovkj1/0bu
r1KtZ9qbxA1htBmTFtlIIel2yIXk+wwafMT+nH1ZqzVo8vDajsPFy5NFjIgVEDZY
KZvorgSDty/LgQ8hprmv9LloexyzaUNElzmh+fnXjJ5hA+XPkDpaA8lOdq9lBuRJ
fZhmMJLCtaRTxEFI96C6ceAk4uml7sApiq42lforwmYnpOsKZz16yEqWp08w7isz
WfZr9P5hUa2r3GqCgEMlc7EC66MoCQn9F6++LS05kcXbIxWaYnGeAXJ9Tsc/rJK6
x5SAaVy0+pFMZFLRI8TkMpoP1dhyblxf6oG+Y+0lLYpay8SJ+6qNHstBbQ7PNyNQ
WqifM2XPSFTXb3Lux94BDvOr8+G1N743EARvx/rhNeN1dIoabVkalfheuYw+c2ZR
ZlmWWfyM6GAR5RRH5zq1sWJF0J+4oDKoC4BX4SPY50wiahoOCNTgEi+WKaeDHfP9
Jhh803RboPCcjNR7yUPS4S2nuCEmLKvb8LHkyVTDNCSFlLXjjKhOaw2KLdOTjv3Q
O8WQnHZcqSFjfrvOBrGyv8ta5nUev5J8MyKzV2MqdWP0tWjBjCh7j0z3HEsmTpyf
ObbVVCJPmS+iL/7JzQqQTJyev+RvPqlDNlPRQqDNBQN9diFz+oXvvax37PK5UDtU
2yrUrz6jE4dKQfkhnItnLK7dyqUGUcG06kPhyApZu3/XGQYSnsjhDXOHJfINqKV4
ysKlc5n5NC9u56tiOPHLobfLVccli5fNXb0hAOUjDXt+jWUNmPXbhWOSTOxHDivd
c2KyUHMmGb7Hi0GdkOKeEtUq65KfKmw9SIUYApavQqtLgOYCb+RNCJ12jXhvPrd6
/Os4ghkwXli2/RRW6s4JT07Nznjgmg/9XOArH9efVIfEwAH1lA2nXaUanijRmmsq
BjG5Agx7TQGm8iqqbIIBAW9M0hsG42xgvkh2JA394+/i20g14J8PDMjB+wk/Kit0
UpzLveqAocdnOc6iujtvoKPvJ2fOtnus6h8tUREcF004IRDh6rf7pcRh7a8G/v9z
AE4psr4Vt+FN8jmPdcigHjMaSzw3Wp5HNT6bkYaJrjVrF+5pyXHQfA+InolrgkF6
Q6miEwu5O4blX8JrQrQkl9PjMtxapUN84gXzZTkP2RHuBmGUOEW726+xLQARY+ow
BOU3KD3PkAF51wn7xT85R3IRRqUgl2RLdHEvg0bfIMftX0ossQ7dv5lPm4a9Cm2Q
wkLL5ArVdw1/RF8XhjACR7dDAuRUHZ8TEOS8tgSRj91c3ix8CYsyZo5zmhgg1fSH
ipiE7DZ1pUzURAIL0TxstlmFnwU1oLoCTh2Q+8CqMxZusKYhmAVMIY9LVb2yyWMG
KeTae+uscRp7+ru5/ETvGYZh0AeeftyspL8kKfGM5PqzM9co2LyLJljM8QqHORsw
kY1iHUZSDXQRWvgtOlg40PdhYACyZwjW9hkM8eBqVRnDzwZ9xzU+WAx2IzE6qg77
mqqGrX0iZRhGLZRzyVbG1E2ij/V4VUDLP+r7HtyQseCVsVv32b50NPg3cJEfabRV
7jM0n/oM10lfve0AkvJ7+4kMp9vKA74zDkCclLpWTZM+WHE8pOUZPJ0mfQ/n7E03
vp3oL5Gm5f7x+TrMo2+t5ITgSoaaveIchZOrK3/B6ukzPg5aY7huG1GCnNQNS6bM
MlJU5U+2AuRpJ09CqxRhgJaYPsuntfTpNWiNE6nlVq54UmG+ovGC8SMH1xzhIiZY
UFK+2T2Oc1Fj0WX6UXDWOSusBlRH072UNTJtLAR56CMn8zLj+R8LAZWKNW75+3j6
yuQ0zAmeRheZIFJ6CRdAKiL3wPeoNOng+9fx2riWp177mnZLFAP5bFRmaStM1Dj2
tZE23tlE65BPQPPPYJbC3RujUG0ZNsEeEePegq1qhFRVpIj9HI77LAFNIcdyG6U6
oF+PSOi/zIaCz4wLJICBvQvt9GmQaD0COpm1jSg2eelH9/bwgZjCvQa1X/5r+ois
EwaDYAB0JJjKJJArqOi+C/oLgitlLpahUPx0LLmajd6eb+F8s/WJuBO13u06ACsa
Z6S0ZCm36zun79ZWL4+r+oXqpieA3n4XUEpXBxSV113NrW6zfZI5UZmG1FC5zOuP
08yy+GOEqsq03tn/UWRsFFB/z+1Bqkr9uDTvYbFj/DlSgZotJRmia4deZyKfwjh7
p68aJVSiP9gff6UdgLhKOxrRp62/kE+LOmI6YK4PmKysEIeM8BJKs6oZRAKRcnuZ
hG269F1TyQt7UPMsjTw7b9AtliAbiffkBWddJE62XmtpX68tG9i4rcTvhYP9DaAA
EP2YN5RRxDCzGvtzQwhrFO6CTUtIDAMWtrMbjncPvVyKMoJrPnc6KODEYLfyBBUP
MpTwLWnKevjmVuLpHIxPrnsViTNdG3RThU8T7xEoSVxTbMLN9frA29S9HDbk6BSM
PHJZWpZaWhnVbV0dJ/jDQB7g1AwF0r3tbBLZNgh3/oiIlWohioWC/RHW2NAVCML0
WLgbgRp0icnmR0XEYRq5S5V+aCW1l3zmZQDpv9Czjxq0NQ878LaItimIz9cObVU+
gtZxeuaiv1mEiPZA68PAs9EM6omwm8gFJzdi1ylZVe6nLrF01DByl1t/hKVdifzR
wyytBlNJe6KSTNKGOCYLpJPRKd2FW+7nC90+OZZOm/EG+KNScH4weieyTWWKZGyf
5hezUH0qNB28BVgYvM6f6oqv4HOO1rsMv3eGmSls/h8ED65+GakV3u04igY0jvdj
54v9BJ4DmKrWIVM/jvUrwjvTKgkfSNgJyKdRPSHnd406ADf4ZFxG+Wk+M5RZLb11
gBZlgFpxiQRaiftsrGLbOrQGIJQZU8mnL+cD1gzLYd455ycM2iaiM5J8bJ9ohLhn
HxD9P6i3AFtdyqckNWNUQZ/7vloUs5Cb0QMnuJMAclLjYl2oyrWnvrYkHZ7ElseL
klVZtY3qaf1ZYBGHgMnBgDZ3AFZwlrrhFm3ltWHORnoFG5aSj5tPCLaBc8OKaUOm
bznygxjy1dCx7OnnMd+NpSeeAlDeYw2QtVNg/hNoRwTY9Rto3RUe3ff7reGGn23e
e2gT7AnDKPkTzIVBWjrASd9VcIj42LTbADbf4Mez+CkSGBCwpXmUFQVkuZ9exyPH
FwrWAQ/qSdEuqzhqYTsLvz8YYk0jvtyQQlLhX0W7Nqp+4SH1vkQ2ydvIF9fKKfOb
Efph9/mNjkovii8SqHExsh43XgG/gMR2CgJls5+gE0DFZMQP3AUTI2zKiSBvYX37
qLY4SArLmptWocetFOveqG6ZycMUI2HbGM9/RWvM6zyC7h8APzc4qlBVphohVnwz
XSLPpLyc8uRgoMa7KnJrTDhdo5+AZEfLd9svUEwZlN0QJrlxDCA2+bAsphWMgeZk
rFDhhhOEK/wrNzSEPIp7Idei8PRK9c+9vI4qc6QQZU2hsueugU5FhCAWyCqZsdWz
rKFartRIO9fQbssfwkpdKd4ZpAu48lsXA+fDd2x0j6n5Oo3ndLZkk0ekHZHMmNYb
VjvanPwr83hXDVbu5pTHKjwsIelxcmO4Or6QBntJxeqHCgn52MgnGOyVK7dRUt0g
7heYqPqT9iye/bGNPGfIn/5B7j3k9ccWMwBr26XFRoa7X8iFrsOVohfBj+uASRKk
D+3qkAsz7JpSvE2y+Mv6OrZlUm+3nsM30FRSWO1+bktNscx/kpyM4VKDNH2mB1DE
M2Sa6T/vxzv/WiVNkuwazwJGN8wwNH8TdUMiydnG9veciKxJ2iU993ST2JfTY0aN
8vGD9DCDIynU1kOY0ERIJ3CVOmnauKdFHjwZ81lrkSsekoNbfY1hXon1LPPsrA8c
e85R2glCxEWCICgGYbWnsQi8yklZnQCIPnS+QsL/12ngZXBvzu2aDWacOFIS7O+/
wpuuKhtjQAcEYlPBFeQG3A3rR7F4k0Zpe+eLntRuo4At0D1zxxnXdX+fuFF2Rum7
LfQnSAYEsyRXB4yP6EGASH/A7nWTr56y+c1c4oJsQCyKU2nZpN2YtBaRoxUpFtin
uXVR8N0fSSPHOEk3wjk0ITvSLMEfpVUS75Gilylpz3qn4QjMGVUywSNoRJ3LBXc0
+C53ew72Uz7f2WaaUuQkGEqJKIciPM6jwJHtdIM357VhejmaY2xNbi0VO4jEftbO
njiQ5aZXMp0AZA+nAuzsoIiVzJGg3UhSdTVsRBlNntgT84If34pnZ7jXOg95BEIB
2hYfsWv8TAlGYb8LUsrwEVnBPpoMxDJM2lMOo2IonoP7yC/ebGcqGjZKOLyoZGXR
29huIf2mRs7cWZUbSkH/TcJMbGI+TMYPW7iKvfXJQo8bki+Y3zHuVYzKBs49ipes
whq3XQT33DVcPuI+i71f0BV5dUBLi7wBZN/6fz8oUxpzN12gdom/Bw3I6bLj+b0k
Sve6tSny1BLenx70YZ7tdWsa9QfKSyMHXDexscCOmXEGBy2OpqWGEBmew6jTja6a
xlqVS2PY1Gvt2LGbFwmzb6eaFTh/Cy9Rt9gXNOPOG8YGqPKzcMQuRWn4TYJkYJB9
N3bvW1b9gjJqvHNKCio92moxMgh0glVt5s5tBaWi1PI3iJDccxHyDKnmHFd1Cu7o
HodWxApw6xepMu9lNBH6ajKzW0/kNkd4speRi9/Tp5R8RPIp2lo3pp5IDRU7taT9
OnmzoYR13PGGlrBmBRciH3QjJa6Pn+EeTxQH4PlobUXhL0sdavJABL1C4gbGGH7j
mqVFFzhdyg9WCgVPkUbLjHl1OIHJd0A4q6YbaMal9j6emV54m/wdqo0kdH2HDx3n
su3IyC5APRaZLwNeSnF38kEHBPBhAoieNGMjBsMPrkMGo4sjXOF5hrTsbtcRC6QO
aPDUafey+rlFgISWjzGlbbYEBgKR21zlUPV66GoTW76G/+Is34asDht9HFGHsatu
Wc/pcMTn2idEXp89VeJwgVTb6LuYirEIXY57ddQPY8EcnsUn5l+mapvgF+/+jKpj
ou+mW2AmkFzM6sUqy/pMSrLzsXrQGNetNFXPyYU3hD7aKgmZw35AHSq77XC6cb1Y
9+pUCGSN8BQ0gGTJlYLDIm7FS7nsavlGr3DKVvN1anGGAXITQa2jrsVkXeZcxgxO
G3r0TIQRgOOYtbAkKo1R+B3XjKCofB5DLm9FQrHip/CmYrRoCbQCF/8pdgg8RQVd
6dVmPljevo7y5xI6cQPvmSjAL3DyH0Y35IA3RrwqwjdCeTWAQBWHnBgk8j4Lde5x
Au0H5/uchICJVO7SOwGTC6I+4CbgjAhtoKVHJEyt5s4eVutvU21UCtclbTOXGaAB
XOz4QlG176MRCcI8DSlYXG62M/Ym1kbqDEO5mb7I877HhUh0mH+8XtnfgsEVKyZv
grAkCLRNyFZKENfM0+VaGs83u/l39/qWgTCZ1CU34uyf7zeW3z1czJvR11UbRrBM
OGTGJ/y/CQ2bFakDiN2Ud8xF0qXD87USB34jrKiwr7YFb1YuJRyhMs13hLkrgpCa
qCwmq1g9D4CTlJPOoEu9s7+nODF7r6m/REVOkdpVrDfH106trylaf9vbKRm3DXAT
4cvkydun+eTvQbz9Zhq2CPYU+2AhXXFInD1xeOSsxVzhoy8/fvcko/8gKnwOh1ps
LRZm9lZ8Nz8kgf8ArxcDDAPPSNxvX/P+3IBQDSjqy28WCaYAaY9bt/blrSLPddNf
qUNlwvquKJAo+tMBICgWw2M/gBpdm1CIiIMrZ/B89cmUWCL8H91f3hWInguUFIyR
6LM52zYEJKzxGubfpoVempgEJYDIIAM4zpLwKC4RKWbuVP73FFQXaCOpaK7VHggZ
lEz8yVdRXSpGczjCFSKKu7Ak9BrYgwAWjl3aEGkGqzN3uH5JbLJBJn2NS4vdep3o
qnmXWzkO5DsJhD0es4+sNZ3LHUhgz4AuYw+XKrOxql/542b03Lrl0zCwIemHAsH4
8RFXe5Dfnsj8fVOppFTQV550SuKLbGUDQbtHV92uBgjbkzAbLrFd7hAQs+XMNmpJ
WYkLFawEK7iqk0XIkmzcjI5OrjwskC33FJJTK2RjYHtQwlz3eZcqtNUnWVvq7Pag
nWyZg5Zkf/8x5fD6yiASeHXFQKMvJeZb/uZN1i6Ed+QnQDzdvOtY9CgRxhk/Ey+r
yJ4xFndsGSJY/uTR3Ej1z/WAI564Jnrs4JhlPujNge8SFWasNKP2rKMkbaEu+tCC
gKtYVWzzmmx2xeFH1BTF0HsB10eqrA/m6xWuBJCedqIMFVWIjj0MqxkjLPyLRMeC
JHU2wzE/HxkK4uSOjdTLq224yxf6Hs4j0pmSB3Zx2X4Q12LYap7YRNibhaZW4CAy
Z01r4NRhvkRzdO75hzE9XKls5aOahbuKlO7y7+v4Hm7cDGW547bgTNdvWWgjoPEH
rUfpE1wMPXXBke0IdoSkqn3YEJGXQBesGD9AptLe3Nw45XLxgPPau3roAnO9SImH
TXsuPAn66s4/HSeiULG6OoaMZ4ovr8emq3S8x9DbNTb4kvisafb5PoevzYEo91/H
mmYERvSE9PHfMgba/MAD0fxPkZXxaaiZ+3Kb2M45qJdwRHEYtCw71aCUZBn3tCs8
lCejEI0B/hz4BFm3secik1MHd7gkDz/w3nviGnRyvzVwfeDDZqGn7hjvv5suQA6I
8qNV55pHYPaCZOj8v6lA3mpbVp/23ijesS9mWU+4MVUEh2NLvZsP8BSM5UoRM1lm
+s3lD1mQq7MFzSj61xqoa0PZjtY15vmQMopMRevATC7oU3TZTcl3i5zlRa91/7yN
E57ruco2colGz+NcGYL+r2+1KTHf/COgw6StU3dSsmNA6NtJaaW4tTwn/L8tslWq
ZyIuTSUJwRoM2qc3O7pqphHXa9Hv2KtpSazy0IW9KQeIYDUPRdugYmqV3k1po1cA
o7qUh7z3IZhaG8WTNv56i9+r2mPbzOcni9SGlonUgCsCIloZCYSZmMBj5S+BaFQp
/Vx9W0iUC4hcFowKnWXCNb4JiAQkLjop9pnn+4HXVqX5tZbRnRCg42EDYpO+HEeN
BJuPE+G7bTVSUQ6E9CG5Da8QfM28T4Botlot5eAMll/Wd1EyAEmT0mTPd10uDpLk
UugETzuu9ohIOBMpeLBzvanZJuZlzxgwLDgxSL1ixEl/z+Kh2gcD93X24zlpD2ui
5ZW5B2+A7qVGckq6byeVf+NTygfVS7XKM1FAZzQsXoPatBpdVqMllYp+FU0x2azq
3K/WSriA2/pCu/IUZ95uFgS2Ld+n5lwWdjLpmDAvECIjwPe9UBTInM0mh+WG4COv
Qo91pO/fwAM1M5n+dGGaufd7T4Wp6yjPZmg18cio3BKhop7T618YSpn7QnMAMPsY
v4zgokgDjokxPm1qRAZo6WVrGRWHiSuyoLBq6rt21Z2E3UCQ6f9VtcpNZ9r7AQid
t4BlI0YXk9vdcc36hp04uE1wfCaIlyEhAUNThE2WXS0K4lSyvOQvtu2cG6wJZ9Gy
A4VjrrmadQINWz3P7PhpZTNf+Qsobv+BPT7EwEcGnftPyam/SLGl0gjIyUBALcF7
XDk7iiWVeGxK2STvEiqsF8hinF90TTChnNMj3PVlyP6YTdiUswLDKoT5J/qGn0Iv
u2UhVQBitT00I3NhCFEiDw7K3Db3qeKAd/D+t8+03WqnbM0f3pWgWG1Mco9zK+cv
J/LwyUKUJFpWdQkS5VKD+Ysacet2q94UH25zRgOKRG73rWNDTn49/v1CTC0yM7of
c2deWT1E0ZGB1bIfuyGuE5TrrNDIU6q4VRbdNu8qpDpqbgakksCaDl3ZmKhzv6Dc
lJwq8KtT9QzamSCTZLK2xdWgyRFuvSxMZpcxlc5H49pBk25jqnbb/vw4FLu/dQV3
UBXQ7LhtEV9Bia9UXWEAuHRSGJpidWbrM4XoQHfRV+CJtIatpXr75nMi9cN8/6ZE
gxXPxA5ciAy4UR0pMbztQuPHy/Ot/HGvSis5XptX5cz6hUrrif9KB6Pl0pcsGEOO
9G9w7dlHH4ew+zjmcxIDbW+nMCOUiu3YMlLYf99zE46iE/Jq18jh92BB12t26U0e
UTRsJNY8H7iAs1FwRfvN4OBih2r6rqRlMmBUPl/NamSOzsI9lLpArrLn+EFXaLlU
kk0CaG172TRD5BPnOdY72HiorW9KHyL6EDpe+vc9Bs2noV6Ssafzs1YSS6ije6Qg
htx0FktDE4zVDU7uFh4TIxY+WxsTR87e8rze0uZ6SIQIfytkYYsjdGiq7tcskVe2
jU/lEIQ4QvcqtKyWzqZT76L8p6g4OsXClUWMR2LrvVKISYl11T1djcWq7Bwk6TYx
IzXUjtTzrDjqWCflUNW87i7u/Tgf+TKxI2IH4p2fPMlgH4T0Jg+FCnIqYm2HEIXr
FbkVj/mos2gSY3Ppy9WhqUDYgwlZTVzXiZUyFAm89gz0Q+mnNaYvjiq9r3HHGOBj
rMbO/llplne9Q+CgoszL6L4n1GZZu1JxjuMNRHm04oU+y1LtPg9BVuI4LDfy1L23
yyQbpt4UkC3WdlHzGlwX+j+Lv2Z51OnS+zVM87vwCdjm66NdF62TU8QwHObNkFcL
fs/O3TJNnYKtCWAKQLEQj2BKA3G5BOOz4SLvDdOPjP7AWtZngI6UOsO0G3Z0JXFA
LODTAqd1OTGkpXV2kGiBm+FJx5CXt9NvN8PMXpDSsA4xo5k3pgXAKfUE++qep3Ps
jacdobiCgBqsYMDxKYqMyuuqCC2y9SN9c1AU0VYhOSKYoeuVLMeiZXWExg4tCnk7
PBbMUAKORqSxcsok8I0wxUDfCwywadze7FT3HenYpjwE8I8tZyOkdhkjt4nRJqJf
uiUL08Wup9XqpxWYZMweioQ9KRvEQVBSXTWnFHQWZbjspsLgCFf+ciS+guLE+O51
nR3bVp8WFLr2uzDMV1xc9nsx8UnHuoN7R/ojm2IrT7L++zP/puwyxEX5lVvpSFZx
LQ/jZmUGCcJTbUi6Yt+yIOORsbYWot1xq30UzXkDgk0CqQr1d7/UggMD0VyyF2vR
2hEmT+xF3JaKPNMioPVcnC8mSbaJCiJQuk9I6oRihRjqHhlG1D/sjzLo8bgV1pi3
KWwnME5UfNlQXxnK/ba0Gjd/+4fewMh77ygZyb3pqkNy64VTzubhfr/q3TPAPJAt
iNng4p/yIVzavjl7kZY1zukhxN46Su1CXgkGhErA1CGMxdunnEplwlLXg3fa7K27
KdKVWEx2A85bU7KiovIpAkWELH/c1r1qa63qtamkOFq3ZsfXb4ftMSicbwc+bha4
I2gqEzxgP6g/MbVEVjyLJ8haAfKPJeYTmrwpCrqdxFdFyuHS0ZRbMYd1/fIf2eo4
pU8heRVZC1Txdq++6gVzaCx1GECF3jmBubIsk1fmrt8hWfxL1U6x8rfkEyczGqCd
he0aLY/4Gc0ToQ84eZyQAbl45hbB9Yda0TwCo5U5JvLIgx0kCdjUWHF61rEAk5id
fSdz5fK8Q5ceETw7zrvrWu7DZZr1brjvbY9rJAldZ5M56RBkmGhTxQmzj0V2mwPI
JVW8FJMftvBe76X/f+Ax/p27axzxIHvrDr7sCxt5P2ArHgAgxXZBTBsN/48JmCMJ
4Scq42oN1wRrxRwofAwtJYqHbHIcyJ19GJjSit3sEi5xVSCNJtBVxT88kKj1gY0j
YNKO1lWCZanNogQGbLhfUT66qB8gNqAKCyQg2QazJCiL8NCRnTDbd9HzGh+eJYn3
8yb3oUscabTEX/0rXuhpN9Dky7LCG/VjajZz8hjQveq73E5j4VJsEvWcKHfphnxc
C4fmMkScqwYTGgF9TU/xwCQlZ669TrWpgqxGhP/t77LUTooomOnS/hB65JuZIg5y
FeBVQx31rY8p3g1DVBAHwXfCTb1MVMqfPmnq70LqhiY2D/Hj/eRLrZ/HUMYIj9Ii
HR+6YpjE1fHuT3nX/teynLzIZqf5iQXvOGkBVrmdgiyA0POtRSEDb4M/qW5vLq/H
eXDcQA6uSn1LzQQGNBNvoRI2vzi/d2yaYk0Y3t4MlMZpsiMQON/KK13f8kfKZEKC
JBR/AgkJAGMXEzyIQ70ctsKxBvcns1PSgdBKs+lcIECYP6rvN4RjBwwSEXouV+tw
tcbQ/08+xYC6mWAtWuf7uLt94l/PCW6ux5kpw2Hkr6spgvoGIJobK9e5p6hptiks
mE6FwYNGxizPMPzlb0Ar92D9E4GOLoWBmDj0e98rjXnlqjUhu0NgdccQS7C5BdEH
FCK1h1Q44D7wYOzS0ZsRq6cxwznVGh81CkFGE7DZJwZ+7olb+BG/j7WtHp2TGyps
azKuOkMGIFcc/EWQQDeJX7JsVCwdsQAph6Vxz0nEWq36+iwnYWGWwXC3xPhXNIW4
foMpUbytQ0ukCqROth8iqYqBhbnECH53pmtTBndORo6JvVJDlXqeZw5gYp3STYvv
3sd0wVleTPpNL3K8LHX3gVehHHJROTQxAZkiTVKg4KenXtaTwrqbOtLaQU7DlHYZ
vujomDe/aU1RVBx/kwAh5UksHk6CAuvypdjFkzclaWUnNBTPzgYgCWK2ZYyoyyBB
wYZ2upvfFJXT8KwfCtDElLTAuwcmUTNqzMAN71sggYznMPe/X6K6uSBnoA73Ftzd
gXtguDu/kuXyC1nLQLNgk1wLqMmQfWvEECXa05L2Avo26yqPkX3dPSdZWib8b86K
9kFsjS9sLiUoMHRgMHuxy/m9ikBrB8Ljie9v5SbXG1pX3pRw3J/lSIT73bcoUUBO
cv9wFd0c+ojKbCiEW/cY6tp1tnFEwLchLIBRKzEf8XH8lR2FzlN3IKQrAXnnWIoi
ukqSfx5ytMel21l0z/eUS90aUCCHyp+qjL9b9EPfh5PvUWCIW+70a62oInWF37IV
UWC584o2WWebCIThvYRFcbcAVswj0SsPZe3syyIaW8oH0m4EqvBT3Kys25KdMw/W
oE1z/rp9l49kYmYy+sXWE4J2IMu3LUv1i3PP8ipf/zjqFec1GeVUdkHrKR7/OpIO
MxsYYJcYgrKaJid59GkAYq38v5VuXEB4/ZSKSfuZQGlTLBx796hV3ViKtia2tnLD
21SRzGCAqSw2PxDsV8n56qLQ/Wk7PbPtof7aoyOrI5UNH2qaXr+tFIcGLR61qqaJ
SQdxJics2Y/8GJz8AV3+kJQtaRktDIdKBQjyXjXXWfY1CvVYvkzBVZKH2V/JxBLi
2GK1Yb86bg9zbUilLNHj9BZh3ZRsIGbDznuejcTbuS89IIVZsHW+iayxMkKmh4IB
/M32LK6ixrsCFTKszpgIN/vNi1zx6Xz1E0VdSmHEDx6Qiz21qqderD0NDDwIfB9X
1nTloagLD5BEXuE7UUBSGIX35U1fX33gpahIWXReKuJGP96HKiQbrK8yEob6Zf80
RPZCDd3pqRX0l+vfOhRCsdFHBpe5xES/8yRFKnOLquUVjVQ/xqxh+P9xIGi16Orf
AHrAnmBjUfm6DwBqtk4hwX1y70MDb75SLVe/BF8jzl5Ibr3mKjgnQGxdvXYZtuAB
Kax4fH15SZJt2mYkJHNAA+U39v1sFdA+WXImJyWLVsE7PTUN4+4grGPBuxgbvx3h
+eMNxiAS2wN8KjErnYk5XJ+ewOBa3Xsp3cB3N/ZQa19TbjBBg14xrEDAOKZI/4ky
+H8RXfasD0nfvq1q6BhOQNeSa4M4whSk5/kWcgubylRSZmQ+ZRRpDEo8h8DhfnV+
MSIqBI7PMP3vkgtBKYSo6uCq7/T4YoSTbjk9Nv/qKGH4nNn6bS14kCTgZdb+gMCj
WLTF0QBYh3sxdm5CVpvShsxEo7PEPY1xPy7rdV3ufWi8h/03Aflq1B6Y6TE5+Uo4
i3QNw0eh+jYyhM73wEt8X1hPwKSNw5bpEcPjPxxEX3CND/NzkPVbMSTpYK0lNmQb
tJr3JyBP7EyLFvlDWM155LDYmJuLUwD8xkrvz2a6Q8Q+hjNYvM24rXjvJ+AxIv2Z
PvCwI2/x1N1ct6SfOZAXGi0tPYF6BYkklDPY7akAhpy/kJZ5nt2NoaFNJhAzmPqI
WvcnI6d0CDoQo1l/hAmHkDRBRv7H0pnDMmrgozhE6WSIf7OsaXzf/XZ1KqkB82Pe
GgZGggeFdhA3WKGPaULPCUFwmTk/a4OrcQjKR+KgfP6ogRrcg7uqXvTwo8Tck+6V
It+Qf1PvYQ55z8aR8TNfFf9cw/otmICzvY3G1V3IzREpH/hkMscr+8riRofcx+Eu
USAQ62EoCFbdrHVuSQN9tyEGmE3IVRR3UCsKiY6mRvPTlxAMpnn1WAEMfvOaim8f
4BPaaNPKS5+iBQd/0vKSv925SC4MgGy5vHgn+FRre4mGVKIKjYwBspF5p7ZfOLZL
x8sqmX41VOth+Dv+GPaX7hzBdo6mfLglDOuglksqkVUCC9TGNKdC2Dt5EBG0j6kT
/CumpylvjNEhSHMeD2q7u5dEpX4ugAZgwDx5GG5Yw8DhEXpACnDGpBTMfi1TrLly
6fwL4jiqQYvznMcFBnlr9oUhWVIys5A0qn6Z2Ora0Aw/gm78riHPmegl9VScKRKc
ADkBN6NxDcPMs7JWJcxvkLDUgpSRDDv5He+ymtw+EijnT6XSt60boFnAcJ7OnR3g
omyC6m+gIH+HXRGiDVbV9bNGXxeDvP/8qEr+0V7whg4kEiiKIDD/cxCULlpwl6NK
QV7s3cbhJoSyETjcVY3DV55AW6sJLIH96p3VR2VO+RTRlvCYaAGtQUiPMQlbjem0
xtrXeXdEf4J2YGI90Dps3do3UyLaAqITePGpmvnWAuM1C+TJ0piIqgFIsiPqso3B
mpAw8lqEF3bBeQtWv3koGbh7x/rnXx85QDYbIYUnBWNhqK7oPC1FWNyEqunPRGQy
69F9WIg2Vxe7dvQBdt7P25E3vUIb67sikpW/r/xAavaPgH0gMqKLi9kPjEgowoXG
SMuQpICHCSNwOI0zW/8eq2n/Ohde/yN6yEwzrqpD2t7m0npPIXjrA516pTi5pv/n
uWoYeP+AeNA8jyRGNvxQ/PuGvCPpbNdrFCb9MOALoYP0w3gC5gcjH+uFuZtYjGGj
NZFRMkieKXKRccSXWTzmuW0U1uazGspC8s+fRFfTPsVvZCIbbcql2QAQi904/Cgk
8BqT1inkEPCjUpOF4C/hmUfuc7FzqGQSWUhEg9Ls1BG0Kx8K/CnWAgNC4W8n2Pdk
pyla8Sw+6eG3O0kqpmpi3f6JmahSNnSgHipEOtNBvReGkgvdBH96tEiKPxBFEofy
0U2oh11W08RgFzL68aAYCRlM7xC46Dt5lJ6S0fpnWYa3v4G8uJi05xKbxtxuRS6K
9jTNipn1lus+L8TCx19IAInaYGl4u6youZ+2dUTMKs3mTnDeAzBa80LKcymuhFFG
SAJgmUiq/Sw9NcJwX8oHHPqu2xyyhC1iWzmvs99JPOOTaeEnbvpbI9DeG4D+16Bo
NNXjdyKc2f7kzsgecsgo5ARaGUPWA9gro/Ny37hzuA6AeDYPWJOFAdeNZa9tv4T4
nbP3fVXW0+I476UjuyTytcCYZw6wLO5II6Q/Sbvk7O+t80PYgnD4vo3il4Z3Thfj
Cdf9tZAG03lTW8gbPR6sP6bhUgZWTznuzdt/yHplLYscQC0SngXpjraVTVBfqIf3
YJ6htYMydl4BBS80revdQz+Ip5MCSKjdhIXnDhWVtarfBdZzvO6zeQMk4ELgcGZy
mqbTXM3GaxFc07SGCyjaiH2nT60Jyoj5BowU6coJjl/+0M3g48qw22sFQQ3muQme
SigNuWqaTFQf5IpZVXtCzmy839gEeu88A+9u5U65ZE1/DMK3AFhrUdMkfe73sLrW
FYAB/1WI4AKzGq0Yx9ysZHsGyfV8USSMZyO4TrbOfzxX5QUaNeMEwpcOcLm2OVx+
5p0BidbrHiXhhLgE0j3n3uJGS3DfHDNBsbRFo1raTs3UHeK29PzPmNLiue0eLkAh
xI7yLOzl5/Xm7QoK5MXnenGe4USSsgkDbz80yTeFbI5RsIpo8qVJluPhszfNRTnM
63Wjlv55BNg6CSdBSni+BGYBXtZpTQ3e1QtebWRsrWWyBz6iHPxsABBRCkBo7K5N
bYGpTVW+Ef50+24wcGiS8d6jn2f6qdfPYax/iNLKKivjNNxHNMdgRmmcP4NMkxfg

//pragma protect end_data_block
//pragma protect digest_block
y9OGA7US87z1KAyTkS38P01Wbsk=
//pragma protect end_digest_block
//pragma protect end_protected
