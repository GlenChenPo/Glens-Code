//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
rs7HEokLv7LuSYeoe99X+DyQYUch7CbFMceiPhY5w3woTncmEi+OjEPQLibmUjJA
98T6fcJXCrfNNHp1+wQRVcttYCxmxjN/fEW4ssIviIsJjCOsQnTnUD8bSxnTZRMA
yhEgswpm8+8jtnE1AfHuEa2O/XjoxApneyKiyOloJV/CyvZ46iesNg==
//pragma protect end_key_block
//pragma protect digest_block
Ex9AyPN17WJbzuTLlVMKaZ/Zc/Q=
//pragma protect end_digest_block
//pragma protect data_block
BhU5ar1/s+ffhYlo8HTqIP1k5EqRiULB+Y55UThaMi/W8qrxVCBTsK6TtcSlThwl
JtwL70Q1CNROh+nVKtwM9/EvkyqGzNXl0v9w25Vyf0J/kku8YTpeMv//t8mtnFo+
j0lc5zpDy8A6JfKrXmLpaNbchw5VyU06atBubzooXoSnDVykdaExSZzitQDR0ZBJ
/Mq5M8uQ3xYQqboIlmYQPYeENNMiLrnZsQdlrZQuh2igzaz6nFFymlHC1ARqoyGi
ff9MqkTvW3Dl9l1Lm79gSMiQqRCRTWMdEPvu9pvNKKeKlUkfqmFtRk+NLDkCdLco
IIrAMPIMcT8yrNJoOcMUJPosYnaI9sUdohGFAgwfUeeou+7K+9WnFIYxmEoOTybF
tSHGv7FHit41eLAIrNDCYh8zP/bksQb+FimBadWdQWZ64Pc1ZwH2Zwo6Wp79Q2d4
uGL52z9qsl/xGauETP7jueEL+kbnsqK/3uLJOn3Vqe5r1KFerK9hGWXVd/S7jidd
+H8NmqHRhX0nf5+LnQmbApGITF3TNi+jCEyk6wLqa+15DiH1P8jLGeiuHvWMwZja
bdO9904ghHD4jP3MuSl4IIfS11ed9WnpNrsdP+cDDl+6KcAq0eC9WZRmiP/xhc90
daBcdgMvMrCl1CbqFhw9Qs63KmJT2K1Fpr8TeILaHhpq/TezPBcSD/gOE9f0ltqw
9xNhn0BrHZKmSulKzvxVZdEMlwmy5Q1SveCD6P7iYHvyA1zWap1I7OwPYgQxTGc9
dgY/1dvKOQanXbKZoDDJqeqk50uWFyd1yh10rMPKbtqnL/N/CkkzVp2O1BpXMt2H
smjeHR3X1pV0NV8KS9VyTP3BhJVeHL8lygLAVF92jm4YZoeMq7mUyULqqivNs4ni
AbahwxOucxE/xRN+yuk5bAZPfjnXNehINQ6jk7ye/6zcTpZj34uV3IUMBV6clNGs
i/7ThrKVhO8KU2zsIkJks0gpXoAgE8WFXagjdeb4qD49ycsrrDaEr6dTckgKU2hH
TzrRIoa9jC+5LDVBCD/sLgWyKmjH7E+lnLQNICv87zWk4yb5oiq9drng4Oz5NcYw
Q6XIqR3JLIRdAj7KGbN4Pm+LNw8bq+BPH2N4xfDqJbZdgglY8BpTRJ3A6unKnsIy
R7V9sPw1Z0BXXyGQuUDmi3vGxRjCnpplee5tPjp6jwA3oB4IIlhRRU9cXBxUb0iB
p1PHxapY7eAy1guzFgrmAQIpn4SsIcfJw9pkc4QzfTFobgc0tkEv7518cp0z3h3M
Z4j+aRpYEn78pNk/TLsxcmF+9jHbi2G8HKWqiJilA+K5wyC7jErCfnpLLffx81Lw
63M9p4Qz7NP9jrs9w7uBv3NcAfnbBYzvMEywzNk756ZlYIqDBt8LeAUuYTlQL+OG
WJSDGUxBuuWGySV6nJAlmi2g0ssCj+1lXDevyVNKkTS/MJMPT3kZDJInSNlibg8F
PU5GI3qYWQQQetPdYFy4w91QjznsQT9UYrWC/mcKHFr4iJGRYnmLzquz/e0TYJ+E
a8bgo69UV8gOkbS6ymWT71e5uKQEqcgp8at8Dei6+AAUMRf5AQT/Fvedz6agJok0
h3p5AZN5GLA1GBayzNLxz93L7MyqmS9SpZFdE4oKaxI/gj17CYLnaRj/5GvOEp/R
trpaJYKebDck7uWNek7RIPgP3tpJxrnCSScfrP2xADYduZdJRblNoz66PMmowpVg
dQOqMO9kcB3Rq9gSsUatGOdPOd5xZPCZGWgCbKhI8cGYXZV7rhYhvtbVhfUR1Syn
0kdNBiYoajKLwMTLu4QTjfBPiurywrajHTCt9cbUKRMeBANMFwh48Nk+CuUsgthY
fMFHGnNf3eHp1871zsPsd+ZxfNVNIDdpvIYs7hEfbo+1uj8zTQuWvZ+Et4S4bYQE
/qopIyDjere1hkerc0KgU3RMFTrEqBQpa7DEuKOdB5jQ3fnhCIuj+W/fv4zkmZ1+
+IOn3hSZxz9SUB5E7c1owpXeuuqNU0TMjhZt+63TMpghNac8ww+6+2ZxUUE7z8MZ
4Dv9N8g5D6O3qkeipJS/dZ+ldc44SEuwGIGTIe5IHq1jfX90KFSv2hSRh5YkhfoJ
baEpte6h1g/LMBQ0guAOpcguWl2tcDpWo5rVmetGw+dK0PU97q22z2FOzspXLNAZ
DR/C1W8Ehdhdulozxzt9UB4b1t94cUef78yH+I+2jy082BQ5keOP++f7cBBAdYnT
5MotD0eQ5K1AMFWZkXh2kY6I2ytwSrlzggXvimefPqqATxaTKeSECG8S4YLLeRoX
jQxYoAUWE836WmbPd12xudAfeYDWyfA+jXWjGzqTgw9J2iCPlqmvdyol6Mam0bfT
UrR/Hs0v+L9mtRY2+m3geHkMQHnpC/0AX586GNXmz9mPolgSP+WTDDWwy2DtetA9
6PS4lVzjg98muHNbHKqtP3BiLcAJVEbUYxMjIy5aYKlKiEufSa+ohAq8kWsvbfWq
uNySdVvkZwjr2XTSYSB7EYqIik1oTZKH0haLtd5Frwk85vmIGTskUcUXThq8mHg1
ku4gdZleBc+MHu95AL7zhoOezTF71gtGGnNB33V1jTlNAQw/Rc5vckSBQ7W+nZfp
syahNkvOOUyzVgr7Tx9GrIXitcSrwL9lvwj3eSmWoRIlGsozh0//uD2hjAvQUSWc
cL1zrFmF9yhVzmnf0vr/OgqbLbimBhmtyf0ZLxrBhG7k7rp0v9z6WSIrd+X9U1m1
aaL1+UR623WiIIAC4ibyTa5Ng6v5mFxUYs7fq4uUJX0oulx4JW+Ea2J02vQ7SZmr
oomARSne0DyGxETzVHZs94OuyluKC3LSck5/2LwOicmQtGciWynTCMjBeheHPHei
7zAz/Yhm6IKYceJmTJFJx4tDha1oirbIhXBUexWRRrjKtofDBZ2+3ovajhEIvM1o
xONlznz+Z/8/497THpobbg7PV02lOsMiCwO7ajWWmAXKO0gT4e32yJFQNJAYF0d/
isB8kIQU9et6jAdJ3BugX88Pad/OPbFnmkpstNSEmvBCippedebq1zJTciT3Y6Ey
nAAcHPbt0OLqL0LuBgwpjv/LjD9BrcrqmqCXEqbGb2HNSl0xSYFNeFGG8+0JgxOu
gUMiHQ3nAZQFb/+jsEU6h7nYKFOzafTiV1RH65jkgX46ob1F/LXnYsscNdNBFoU0
0XHzAiwfdRmDWyGc9M0zTFoQVmGGUgSeYz9NtSscopo19yL6IoV6SpNstem8fVPk
urP6yqJzukA/dkvm08xve/s1B/E6J7qhdiOj1VFSF1H/H1NsifTscyKWEduni7eb
DNHI6/LoKME9dXviAovOX3Ui8XOaVFDPsT/gZBgbINKcSnbqzqBf6L8ozqm43G9F
u4exoIrHpBTcETgjX+bAOQWMgwuBZ+c/XR3wm0zPJiYFh6lM9BH6T/HXvn/7vpuY
EzwTCQcqHiWLlintI7R4/NtKBiycFJJBFom2JB9tF+OelxTa2s3LYoO2EmuXiCtz
NCmDrcR5+y4qaM0NZCRf2yQB05yTwt0n1XcGsdvZLHolecFbRiAwpnY5sQkel3V7
qDIqaeCHlOS76sc8JS0frGUQWynOxX/9pIwO7fOgLXjH1M/MBLafPy85xqHwsVzZ
0Y2qb8PH5OmHkeTVD+PcN34jva3qvH701hZDWGNbC4aF7Eeu7r9879X4ftkiVH0+
adlu4EWJRP9XU3dAd1Dy4Ws3nLxsAOQfa1AUaovx9OUx/mqsUfFhxya5e88KchkF
q5aXdmvmXfF+fu2clbNer59hrVkoGgEm0xaaoOy+K/89gz98E7cCg70EgMlLEo6b
1ekSdsVOVjd0aJQ3ui2vk5LFTrVmE4n4kkt4IJ+wlbOkxqA2FDwnP2yvM/t9SGdc
KrFCnJzuJKIfhqgagDP8c7Ash1xx80Jcyarp6ULDDuwdKpFXDfDbHhEjhhpEg9v2
MjpCqzpZ13roJQ1O/MRD7kUBtAKRm4G7VjdOrcgSQgUYtgTRB2IFVihJRwUyayP3
EJMOFpw+w8E+jEI30ygpT6upBbfPh9eLDdGIrXR07iciuEVg/IPUiydKg1qsfgDx
Sa891IpG0vY172wjzm1ei4uPhiUlWZv0Ab3qzVOsQ9eN7Km4yHNqF5iSbK4GUCXj
c5LpszGXolztXmQ2b784WPea2fZ/eSzPhQcY+PDw8RtgIkiLUg3XKETZxGR2AbH4
d+l5i8sMWNQZ3lwRz4wvjSgINBX6oB5kQckfa2wTZPvuyOkpzEmuoynPf8CQnn7o
huoOGQLU2D8+wXKwQXLJ5sPG1aVJ3ZItl2W4xCE1NdqyTAKSLI5n2QPZ7Wr90BZV
XLCRcM5BRcHiQAiRi6FhLM9IF9nFGsBNCn6WBrUyBWqxPSVlEE8umgtO/kiLowK7
kPKiwk887J4yUGtzhUoGh1vTiKOPk0/YIMkqpJQB9Lrh0oqctBrWrj8c8q4zc3gQ
Cz3LFZ4GFV8roJWOdwiwMKEmeRP0AeBZX6k2e6LjUWvml9xSG5vA6H0sktuLlY18
LJyXC8IxwqyGeUY3Zg6JxXLYL5efnZEmy+JdZYsoBlYKhfxLIgC5GQGmwhXwkswo
s8MEBhoBpGTeQoidXNjESnzrTDq5ngxBKlCroVko0e2mt9ozVNp8dLcgBBBHde7P
VdOwa3G/uRx2Se2vdpz3Uh6f1I+SpFF0CA8qMqvEfhGRRXU59CMv5g3meHHAJUmI
XdWkyzdVHZkDfVXHyF6M2hoiEBRKU9swUGEgOQzq6oOehrKhnZov26U5n8B2sKA2
cbeoS5qj5pV7J2JfogppR+t6Eyx6SE8VbWjx+E5USy8VH+3xJRbyHGB+mQfD2dE1
fnZVY3ikzQCQXA0CBqcnOPhmrt/+QGX1jHtYaXrZl964R4I+9hyRBqgcBm1duTha
lXdooGohdKW3kZ9tzHx7od+JaDjOIigk44qkbintcPjKNuly89qWEZbkLEuJBBM7
pnOpCFm7xqDCsrmO8UvasNCacBD300raxODLUjycayN2q1EybnlWWoH7GYopC9mT
4r9v/AaVYW2U34yZmPFMjBMJx1n8HB8cEHgEoZbS+DZJmLJBk99CMr4yiHpConJm
jWzMrf5rFZLONWsET+8UMtcv4p9eK/NSSmAvbKv1Vt/47BWVdV5Rp9zwxGdkpO97
8QnvnPAQ/Ca0k1dul4n5My2hwvnzbR+J4M6J5CqDYdBja/V1aehUmw0bHnmEplsy
w/HvVsm/QoSdvnQ7OmkKa1ROZCTraqKng6qYpvlAHqlUpGnJjoNbdFRu/8mUqd+R
un1JJWVKAM6UgR65el0s9R49FeucIoZ0nbY2A1ptYhawH6ezhlPZ+mVvbckiAU5q
rm0lSn3+ii7GyjyZvq1y5oUX/Dkp92S1iAJvOsX6rM4L/hjPI3wA+0kaHTK8lqFF
7Rchb6Cp/vXAWNWx9YuzX8J+FnO03dW8MvxdxNcOkwy58wEGrW85w0YBm5DTqdx/
exM7P5SJpr0/lyo8OD2OZaIbI2ZwKl3tMpy2Y1j1SHaxXRJrfshRVwJcLPaE4y6S
fcDL69eHQx8l/2ZohrpFpA+VKtjH1Np5PTBJjo0WuV2X5UJ6oTP1eeLY4frq5ytJ
BaBxWZlJIrkhdcIq9Q4vlMNdO4ESNYLhhW2qP4/cEEt5LF1dsknpUlfj58AQpQhw
1fpaKyOO+L5Ah9++9BNYd+ERxJh8CcIvpkiRk8EYeGXFrEJh4XLKZoy+eCid2VWa
aYxyv742Ndlz0VYGXKdhzz5cFsSDN64lk8aFxAreS6FE6Sv95Yfi0u/EaF8NIg1p
avG3jmYLsVTdBkF5vGATPtxMLvHfsp4mRNe2dKicdqUEjejtnsC/QBAEGJ+ud3BC
ay8hswrwzkVh3QW1XC3gOhBEaAdHGjR0UFwRTFZitTVpOQ1C/s51W+n4WMcrRyEg
1OmUz8FNozoX0qXfnebyGbwyauE8Ijmy/lDyM1ijtVcrtXN+fJ9lPxpr1ORUTeVA
bv3/wP8Vm0ZShpjiSdXMKHN295E+1fue9JUCJO2gKFlukhFzkBrE7ZnAidsoyvXS
9zrEdVKWOCtX6XwVyF0HIpCW2ZLFCGCGiEXP/Q9BZhPJAin2zRhajD0yAiRQrwkF
PCcHm3jqJRiekbPvniEFtTFfqSTillyu76Gnc0FxLddKkZPZRWCnk0tDeoysNmpN
mj9UggNw/sMfQU9pY8AfFUsagjncdYao8j+l+zxfU1LiWgRgUq9Px7q1xusz11SD
FFB/C0YjPtSyj7A0acwvWCIYdjuqB+QHVToXQukHnc7Efx7IgFzkypjg5NkX/BOe
5RAjgtPmFVz7XDzX3wFDecljqPPrzVnISAJwP3lAVTr8vKCOqnvKprS4DTkfrR4T
Z67VkR10kwd2Y9BDRd16RavSAUyvSzcswwAwhkORmacWa6gjyxvxZrczLx/hDTDW
72AoI5zsBy0S1IEHvPdquX2T5bC3InQ9EaM1w6jndpSzdIK9FEZGHvyFFjSJWobn
z9qZ/hl2MBMtIgKgfIUVeqXfVMFsivGo5pKLrF8TARvcGQRn24kTC6WhpREgDNJ/
NRBI/1nVrKfRfgBiY0wTg91vSpRiFUdRGduP0vXC8AbFQLZSagmapjX24FkuLZff
ynEDPELldjLc0iBLTlOLz4zbqg6pc5kSvRy/tC1Kms0HiVYY7QbgwAQGrbxtTuJY
kAWZUCzn5EpZgW/+h5uKvElLkb0O9Du27x9WjpL3Ibwi1LSFxm5RWWbR4AeEoy41
94kW3LFWDPCLq3u2E3FqLQu4kJwJFlUKp/BNhfhV9CyStLzomvKC9UE1wSMPitBW
A0JCgSNKJU0ZLUS6rMmjp7czR9HlnJoH6r8FZbUS0EO+Kdt0IMM8ihlBOjX8+SYI
JD26nN0a1qNx0mAyE+eY/ZuJsYt8xSH+x8u/YBeIrb8CjNFFlACax7P4ArI/mrZ/
2qbGh3Y7xX537Ypvw9otLx2/kjju6slCUB22k46FTXV0zSULsH5lf8QCCIkHBrM5
PeKGSzdGTMdzse2V9tQmyC2Csb/g3RE+PXZQtjQvJ46zdYW3dA0T7bVq9fcV88Nn
UyCFfCx5j6Qawrmpu0hKyymDth+FPoOuefVkjaAKE7uc6g/C6ufWWPv/2G8mwHDC
SLOLzlPRlBNWHDlzHDpSZTWQ42xnp/JETLe1b/IacTj81i9dWtXkuZyVEQyg7bNe
jA6Tm0LpS10kCaRhdhL/BcoduThhrItOXE0myfaNvdWg/cMmsNa0wNilFF9Ts1DJ
iqR2gEV5fGj0UJTVE+gQya4I4XlFeFbzLEjFeCkKG5j2jM7VBrmwAY2DsGDkcXTZ
hjGt7GIBUGARrz2lgyYa/EjoNo3TEn8ZAIKcaOi6bcc1bFxFpVzkhjZuRTK97f8d
y2ffSedpgKlW0OZTOek8KgFvD5q04tlOIE15Qq/o2evEaXfA2oeH35XZtG/esB7k
4VwFyctFPqDaHTAIYGtW+bVmbYHcCRuUpRmCwbV9w+DTN3GUSMAGMoUmC4BluMFI
IgJP1fwcceXqMpeolEuXzaZz7BtwlldKumHK52CiOqH1ZemZ+t49oMz5eX0iV7xP
/mp7SQoy0s8rJTvooTVMY5oHJntlAMeaym03VPzJil8A3P2W/8sKUC92acDWEWha
DpLscDNZtve3lhXjbN1vhJrBkkVlJ2qkEYcvqBjviDuIEWwcDbhVVseAgVS3hEdq
PPVwtM4+yNixMOEuQ4HAI16esKF2jBbdNVROySz3kGEr/k5Fy1kcFqx2kDtfIuxp
bLlm08P2acJNe+a0Jj+RDUk3YG/ML+C3SILAubRNtSZ0q+tRcAIBA2dwLgV72R9g
GgCQ5kRdo3J7uspQkEIdi19+7VsRstj4BV+zWeyKEhkEGGxGluLi32DCXxdtljz8
32YDbF4AXvODZUfpDl413bg4fWPAzDa3Tu7Q2DIpic9JDPr8IkPPf3UYlduybD0V
Z1QWv85EjwRAadwfWDTWfogTD8fpkPhuRlOY15mvLNZDaklXjs0FQQy2ieXoC1xw
nvXHTHquc6z8jSjhDKnLst7rVnYHTkgTeVCW3On9O4Vh9cjG/cTO08boxgx5Lkqt
YmxEmYhwxOVeXx9uxyMbZktnoz7TJRYjYY5KGmTekycfIVXgwJpwFRJicGo3WMPh
8JEsuKMofCIAkgW7anrSvBzmxbhhTcDBZ4/G6aTd/7j4yH3xJxEfPi9m7FTVuU/+
XeSb0GGTKAMh92DfU5OPfYlRtuTvsvkRcy4P2XMzQdo55kdimUKtA+sRB1fP3y1n
3ud61NtbBMLxhP6e4dSDeXmyY8B/Tz3b2lHijfg+4RFvYnp94VOtMJd5wImp+G+2
/qeoYcbplB628+OmEqlPdFVCrrtRQYcymYKaSNlNnW8dFfniC3jEzxk5jdOI29Cw
qdg3fRBMmmZAA5OXsilgLcllEpG1Fp5lfKwGbOcuNjDwHIYy69enZKDycpUyOFt8
6OwDTnSa5MtqUbZTg59F1Vo58vQOuIQ+nwUGZyVaTouwOl6rkRK0oDqp6oupNY+f
98msxL8SPXePwuUQG3Y2h0lXUxJVf+842W4uvGjUI3vL6Udl4Kd/q/kv1vxYYVOz
zr94JAGCm0yXZg4YIeD+etpYAufaHsNANtRs+sBYvpd0MII6LRy9Q30vUUs1dLj7
9zW9ksW8kwpfRBu4y81po4qpTXn5kqlFUVIKbS4V3VMg9RCMtixGX5651ACCZ6n5
8Wnr/A+9WVV1PoudnMTr9oGVMDFO94EPGizvWDdW4nsTbNp7GReJccTBo0gyhcP8
h4xAMQjAkdp7hyjR7Zpt9zRpY8X54B1HO4jhKF131UuE9N+i9ytRdR9jfzvTwJC3
vj2oUuzqxEKrSxeGdL8Rk98HQ+Zu0vcAsR5SFIUuXOV85fnN9Itf1D1tmrJnitTj
/d0eVEx4bXuaNKvNUqHH0xQaKhV94XPPxqE+nXLsT1oRF8QAwl+KibT+gPhzikAt
twu+x4TiNJ0ZUL5c9pCQZI3okpjwjLrc7JHmJJmR4mfKeMKrTHt3oB1qc8R5GN+h
LguPPYfp05zTXwQv4//o40IrVSvlZFqBQ2Qd51XTyJhaK6WkAI2AMzkPiMqivYkR
G3IGkEKiq2wP7aSR/X63P35mn8juJeogvO472dT2M3t7w7br/6G0NfSVOeFjEQ3R
7HRa+r9X+ztUFx705sDBZP3j9X5GcKJEljXBq1j4Q8Y+cnPnZ8L/oAOgnx201p/v
xQ4EYwV3dp8iGyW8cVY7od6byQqYIqTYIPVA9ShkX+GuplD/E3fXqBb4TtAXq9Rq
VU/T0eDPf5Jsi3qrrcjOqI6dYNq/nTpzW57FkcxOS25whPE9BrRM1gIbf4ifHy5j
8oB71OVycymyrpXDfZXEXKNdaRTDz+mXgYYO65ZtksojrKuWqxr802vV0v0LTDkO
FYdrCbwMUaIApbUXJ2aOWkOODu57BnQhQEYCDeoHk4z4swGnY8p25xJWqlC3LGQ4
NqEm9a6RRyT8korXgmq3njMCkTMJNk33ACNt4ExXscYDXjvI57lSZPGRcf2hQJ4x
0554872F1P4s/XJVeyYJPX7oZ6E8QSdLcXfqwGPNotgDLZtdLmGt+3RjORXROvLH
D2Wol0D12Nv0PVwanhKX8uZfhkk/O9bideJytJnvCoWcGE2lWHO5DkhPm0mtVYsL
h6oZjEQzo03Vk6HQ9dwPgOP/4/w/psTrshf3/mXdQtQ6UF/S7xR0UAwVE7RFnIY/
1uWvhaYFgEJnCwjiBxGzz4aca5aBj3DnwL4xR62qBW0UoTPAQul0VvahILaHExRP
NqMsUIWYqRi2gPe6udh1TnZqKOv/RjLC0X9l01Xr6DV056VjhzLPB7KieJ8YEfzh
h70E49SUXpIydGyBR7XhUrdd+QiDUoIP9e9N4RLO6dG+Xx7dWm9IerHQVAbjLP+k
Yd7v2vsCTmlJ1xuw7r23tt9LZnDqZ+6Fyqmj02mf9bAZkbX4sFGxor5TOPZGs36g
KZc1eFKV5c4+3XyBysOfPkb2GZYedQQ75K9jlmVB1bpyeXZ4afCUJqEbECoqetYe
m7KvK1ihF+2lWOJ9MXecvhF8K4uDRCydzgq19f58dEHCCaIQzyuf59GU4GT0XvhI
bTPU4qVzVKeCo7ykikmX9qR9BEp7VdrkygNFEYBEjCpWe4SxhRJX2xUiZzgE6BYU
lPnWaVlPur3vjuCF+y1hvjypd9t3jtMuKPfio9EHf1b0QZPqp7wCaDMvI+kLisTb
OXwpI4I/r/cjdfGOnWvRMA5EWWLg9Fi4QIWR0yWd6QN3dPhEGckKStaAUcInlIH3
c8ASNxFWScjRhMp6hccISy4V2x5g/tWXNXftyse2WKStPIEOvbB1cjYoKW16CZeF
aZmAqiLcJG6ZZ5+GozhmlMBU57SYQUoXhuExLwOi4z5MJ+HLrl4xIqUFI/Vb9zx2
16BNZJJT89sdKY8f1jUvyEK/7BDxFwixb7PdIWDgQgpFvioenalKSJ9lS23+ocdw
NMpeQTrS2QeSNJV6ejEX+oH3qE6h4gKVUI51RZlShwRNu6No3xl+puCcKgl7ijvb
bCe+/91UdN2a1BkaCnhx37LMjBnBnO4VAJ6fNHYeihzuW+PCIJKDJo6BeUsj9hnY
rwfID11kaNP7de5YvD9UnyC5zOqZ7DbzamUvIfQ5rqnrVZ8FGCaLi18eAShWSjqF
8xryshkRJAt71G10PVxClXYEDr35o2Eb/Zo0MR81KqXU7apwyGrD2F654gvfWOmu
XZO5sJCdekMt7m/n+lcCRrspGcRfj75H3/XedJLG4J52p5+t+nUxWYm9pt37l5D+
RtXaicX/Pu1dNyZXozun1O3iSmGoHpnf6eY6UhUQfKitPmK/O8vShCKQANk9bNq5
BxXnaBE7YWdl+VdP2n/3Ek2gUC55UKPmI0+8Z7c/mQDIbEqpZPNdSjSI0pINQ6cK
5sycQ4NFyM6w80973lNl8LRUJgIRaMV5Wr0G2SMY1+FSGpVmTaqtxInnYKIgKMYp
tc2jJipy/GckFKS6XFyLDHpWln0Hr7VvgJlMB5bgQejnvZL8JT/PzmKVfwdumtEj
HfVOlp/mOl3/ZFIMDiNhIxPvmD00vG+OmJ6Mr5PZlp5Yb7d/7AfI1bIliQ+Wv038
lgdmjfiN+JmYubEhVUSFaIv9G9T0g46X69P5y+XUu7caTeWWS4zZxS49bQce8jRV
WtlcovZP9lNbshj0SFo2d0v3cfqQkwoECNMB4AigG6sGjO5eacq1OmLCMeVdHZMA
RebB+SfGZvXvb+V+tes9ogMPC25rYVnH/5hBP8lQ+ZzACnEkQZQ931EgkElMo2Rt
RKAScB/tFfF2JyzWdPdzNNCcMLcfaGm2J3B/efQiqCg8l+plycfLpL87G2pU6//5
XCT5JE1S21+mtVOlFDX0Mjbonx7nly5MscjFyGzvfTc2vPxP8TCmsnj3c5EbMOGE
lFeVqBBCYB3+5ySUlDrzwbErUboS/P/5sqhFmLzjmDn1d1dbXPRabce+NJFIfMzX
eKDGpx947jQwWZXuzibrR+ZfivYfZB93YzwXPDPZYZcVd593d9Lr0g9ydi5hwK3l
Hhia82kJzypSx+AUnb25X7jVa6Rk8QPR6BedKsUtG/9klZHCK3sNwPAZoGu7Anji
Gti/g78ENtWDqzW59yDkNX5UtN5aAxZc9+eoot0PV71JZx1uo5k9ZMr9lP2FxX6g
UQjgY9plBwvB+zCkaL4LVJmwvHE6EObTH52AI3YUuNqSAQrocd+LagYTZYytTg+F
lTTiD0kCNKeh0NU90XTLhSav7pFAt9spXmq1DYHw0QUOpopMy2JJOJ1WG7xi6bIM
kOgBqITXITAtbBvv3Oz15GbMpAnUR6dLu5p+tPG/e+vKkRB5D9InGfcLQUYG4Fcy
EfqKoW3xcinSEkpAvDjWfqoLmXDULbVWgUEl3gYn1yqUA0PNxPpOzJx5cUdlmkuk
90sjz0aUOzX0J5B074uAaEm0qPnsddWVjrbwiOTJr/cPZ8lKrCVFvPqAS5SxDyU1
Epx/2/5XaGN7/dmKxaMkFVmMHZ61pqBO0mf4g1qMQCZnK4I9MPc6BCl/JBbPt09w
yGQ3WNXAxCfcduSiYfUrK7wd1fCI6+B0AEuYNvqZy6gbRwa6FVqmNiowyTrf+eYW
2lxFbY4hkSY8UiZDweORK+gnDG/ES08Z9TMYxrX3aBRC/0rG1gHwvzZF26TTSIwT
83sAFghTFV/enzQFYri4fFkvteIgUTFLtyrEJasA32VkfmfeLPNsvTU8eroSKpFk
H73VS30TlNpLsACC000/15Rn1jUHTzjeya/Dd9R8kOmcsc1NNSFAE8Nj369Kz9wA
04Yh0E7hWxILiYz8FoPSW8NvHVGojH9wvH8eDqN04uQw4oM/he0yheFR+cNZM8qZ
zolAfYszUI4tOmcwDDzc4lokaOBdPzxJ/uINKI6ndGMZL+Ta7l9EonNK6BYbnHGV
3CVDBsrI9SzZmSJzxdCnSBqQNuz8K5/bzLxpatQjK+dl9aTzjHC2thnnIwxwPSag
1Lxbgu4v9apoozZMM3UfZgqQkR9gISMYlfC04SUpF4als1EWD9GIwR0ryMH3ou3j
jwvLUAQCrscd3aJbikzY4jGhUFijap5cltVlbnPUTkVW7LEM/Jv2Xb8xVeIls97c
ApTvFu/wyAZjX+VLoH2kFKH4IlQGY6jc40oYQnGs8q0plBuSN8o99WXaiqb6vJ3K
JaRY9eV0p/r7F5iRDXAwShjRQQ5jUch4fSPfU/V+dWUc9czncwxdWDNO5wYr8Wkm
Wtam800gbd1W1s+Bkir8kYxhMYLtOQ/mAh3U5a9YujgVwlzzwjES+k4lkPiIN/bt
HjngsgPh355EgCB35+B0VfDvB2QviDQ1Vr+vpBezUb04t2yhthneDnXscZaEuugB
wy7D7g8mGXx13WYC9/tsdHvO79SDbxuUQ/8SA3x4p/DfuuK2NWkIFcPxlQo57tdd
Yob/4v+e2QvE0NVHcFPFpLv4yomfYeiT8hlL58zIBjVZfvO/6uji05QbRXvoHNYU
9yWSeUFD8aoUglaatn2lAAczuhEGdfFPZxmaNSj992UBqsueXFi4RFZdkCJ4WxCX
LVrIko60Uzn2O3IvzOVRk72Q/0dQ3wc6LuW2ia6/U7r8t1LWgM7nu1v4hk5yqkz4
WjszfDCklH4zzqjSOwrtLOnpUr2h3lcRvWkBX6vyWzB5cHvgYbutQGaNn/8bLQ+e
AYV8y5qMUHZrbeB5qcnX9ghqaVhSUiSPf40fEgvi88IY1ZCHEACKo688IPWfc2y9
o52en2Ap+rbZSeU6nLMsmdSWiHOCIE0HQh9l7gvpxGfqCGtmWhkJDulW7wn3o8v9
YX72NWQfp3/CAdowUGb/Uj9TZOl11wH3Ve3QcBkOFlEQEs9xAWM73dHYTdOgRjTH
VK/obtnKyT4EuX/LAXvkwx/Uu2xolWLroBkSqkCC0ontxYN5xx0LwKFpZfh3WO+2
Y4PQBblKu3EA4UT32HpEroFoaOlhle24RzmClLxvgGjsaqJkVvuSxrb07EihxmwX
mCjCjmZrdkdgBla1jl29yxXbpJh3D/4pTGxmPduGBJLf0w7Y8DmxtLohyd/0mfUD
qIb93e2VhUsxSQ87D4QV26lETOupKIw5/DlwCAnbe7qZvY4aafP78KegGyCqYlOc
SNzSFmzpT+xrm22uu6OJLX5TJ81iLqsr9w+sTXfYGRNH294gZYiI4WIKZA6veEcN
We5IPlRvEOC2kOZQ/SeHexMNK9oZzTKa4H9FLMbPmEqt9VkdUPHIUo0JZtBtPMVN
o5rjXSUduxJPb2kwd+QNS69fV9NLeKk9tmCAdeEQt1jHaGaMRPcN42rCIvbaqQZt
XqYZODQdSwA4oTCZoGf29wwH0F+HZCgQxvzc90TkMi2Z1WRt1kvQUFcN3bSgmU4P
Uy+fTgWRDQNADFXnTFa+o71SUO7b5ZP75A00DE3tKKa9ulGucjtACDLUljJw0ufz
jwJCG8iztMHRR+iagEBauK1W5NkN1+8CTrQgrqNXUJry/erPaO+6wW8K3wolIvaA
yuBA+vDbKHGkoi94Lyuh4I7TriPD3VQ0HguUbQIHvd+dHWrWLbki5Z+TnQLJDQE4
gyGbEviL9/RgFE5pozRyq0Hz7ab24/6TN3jOi+/mM6its+mw/0U76uvsoCgS0DWn
cHiEValgTGfaHu528ExnmUaLpGj8mWlYQyn3QlqnRREB/JGwl48Qho9bOqtyiRgD
V6/gAwIkOAPPJ2lvhH/NJS4ytIDk5v7zMuSUkMem/7+I/KgEk7FpLBNGutz6vlJm
GMDmgMn0hPhftj4n4UBxrDXr6qB35eQ8DTXZp3uOuSvnD6o8k8i6E7n/BMt4RdkW
ArqCgYuHSXHTIjTb4Has7UR7q3nOd1xj2LuP1mawgdpbxGmtrGGxatgDinoMS4CI
HvlkQhqmpdGb+iVLpGZ+1eNOOj+c8/PrZSqpxfLgd23hBsxGTRC1gkCL/V0k+ObC
3J05B2SVKursC84VlOjNLb4DrduBY8EbO9d/UnKTaq79SNXjyd0Rq6gCgMskmlid
R32WYkICgKrMbj3NEHg60HRJYUPHnT9lIuCBAFz1bTSZzAAaEAVvu572sAOX+Wlg
g46pYPnWL9WuHBLmcNfiBCtg448JSoYYSxtXzIKLyoSHdSNd6mQQT3SQ80aSOXze
atggKrEp3HpTXE4z27/s4FlyL+MuMCS53h6Hp8yzb3dE+kB4LknDxBIUym3d7mJ5
GifdlHMCqM4I7rIDmXvwJzJhH+JhZtsG2G3IMyLRJywGYCq9pDPckaWx/TPuAZuR
dfl5se/Nst0DVsKjKoeNt/lJEYcE9L9BYCNL5fbPVJ5kAXjyTyyDcEiyZhWyBEop
QIrdJsxqnHWUWoywDLkzQ4PRHzD1Trba5nDVBEDKURX0uZGXbxX9VF/RrZfKUrUe
BVufEsl0YF3gJDbAdkZygxpOSOQkhJExE5QZS+304CF1mcnXm65FKqdYebSilmR8
kz2soumy0BO/myxAxQWXICRKxD+NYwKYgS0Ng1rt/EZYcX2H4Kqmyz7Egw/uXDrG
1vJfzl5tP120t+iA6OCF5Kq2gXcf/MEMceZe/dUhRLhTtzRmbDrz4dL4KWD48ATN
+9LB5Xnr1GHZYa4Pr11f9j0e+Ps211SEgrLxHuU2C/VgeHBq7ZtsgAF1r8UKx458
MHJwiKcs/BZgHaVUdq1jmbmxb933NcpAmcEyi6e0BLC8wc7d+vqLQln3nXI377P4
zL1MoNKx6q/KjkWx8oU/4TgAvtOFgetrbGf9gTR+5gXHrZikzaHJYum0fnKEEDdk
+FP3xwZVqm3+A35WjyO1L8/vBdCVXPgt8UYNT/K9M1KoLGIyUDbP1yXnBWs0t785
OudYoq2dklAWadp5LLs37IFIetpC3yWQf3DqgK1gIdCtBK7Cj0384P4wTxBrYrjH
k6ePvPJGPSMIPXzzhvO8ZJlWbDWPU41LKFaRcKCkwpEjZ3sPsG07nD+NnQCD0Btm
OOsawsRx7g2344Glx5C5dOg9zegRKJssb/MVOa+fZ4ufqM9ehCWBh7fgVyObXAnN
M2hAx2zWrafeNmd3L4UdDLR37+3/zvpNrObbQrgxj5A34N6t2xA/lKQ3WxR/OIrM
AC2cQUgDWrhRTRpLLMjU1OJSerZvuZLo+UOhH7eMH6PbPEYGpWNWN4oZrzEuWV4x
CEZoMHyS+gOmG0O2AcqZsi/Ysbf6ryRpfWXIrK5qaEOWYsRi9t5Zi1o1Y/fqD54M
Qs1W2Gct9J/ZeNwK2DAZB66wXtb5XVaIybUiXVbekzDa5eYLmbFtI7WCW22FXqCI
bEeVlFQBiMmuxmcRnXXNoYA11qDMC4gXBuctEtLik6PigtfPrBgp53xPXfycjFDt
SCq9tKZ32rrAv0gyXo/tMQ8W13UJEufplJM0dsMm+r0bTCC8EWQ/9OKwQOM3i81r
A3T+fVMEIOOSaqx6p3rUODkV2nwjrnLPjGaO8oTMdNO69eemyg8qPq+K161A5Z2U
sJlhn5MSi6ei5lr2Yn8SfYz6tiyjW6mqr5XRYopaghK8/cO7ML37AX9rMhQFb/j+
rqDRSMt0AADg8b1yJGXLt0Ga720RMCIHkXA6XcicfBA2G+qw+HxA6uGI+qFICk+Z
MKoDo6ZNDCyYKJCJIimuqgjUrUF5B6lh5zFKjVhamlLcTTZZEzUsSNWH1ClVF8Io
7ddcvIlq5rGi/SecEwrjNqN2Ul9tgawR4Ie9uW0iIR8veTGT91X0hFeRuQxa3v2a
56yStKbh1j2LsYdht/ilh/IU7ppKCvkt7vY+jrq+wP7R9Gtv4ij46Uc1omLMeT9E
pAKA8IHX/ViNyQMFvU0k9zEm+9ASSsnoC8Nt4JPdvGTNr6zHxVQ/HijLjPZYkZqg
/F6wJ5ZE2gDGGJU6XGdcUaxjhMl0X7hnD4Ynsv2mtMEnbzwb8OtXxwVAGhi12887
oNcmu5q6RkzatTTVVv6qgFcx6ZtuV+iVlasaswhBdf9gQ3qBSAI6WFILE4wrHx59
RQmV+3mqDHIHY3F+CMgQ1NwvFZZ7ol/MKZPkRoxqGECn9ADDtaD0tcExAJkj1OPs
0XZ0EGBqPSydb3OzDb+PdDD+/juhbd12OcyqMF3a6MVVNF6ngvcy0KlaeWDr390r
p9MU6td3pCxx/hfvQG7DpCcAMTDhVMbb5Q32lhxeykom/u2imVTcbf2qWx5VHiNL
s36dbDUvnwrLLh2+GwnBuPBFSQhwySfEdRWO6eYQBhZtBWecNPCmxctG/T00Yhtz
dRfKRAyd7xkH3oMaaiPdrp5QpKHjTTno0P2k9Jp9NgFIz+0/aPi9XlSINPOyNM/U
YfiFJoFge2vL34HLTb7PVnuLMmoTLOjYaCQTH6TXL/EjaIK4wPtCNQsQZ2h1rorO
XYh6e/yu8oC+9qJ/lqdbc4JjwXbl51EXsvda6Ou+YSLrbAYPho3C+iwkQBJAJZTp
UCnXusv8lsm0kRfRlKiLaprMLTM6QguZH+tL/5AeMnDxnCXyGtEsud+KwR/9Fx4b
IMtmCddRp4WPIgr4nAjtX7xLW+7/tz4oJ9GxtcJ9jesVSZapv9exmzO+g8iX5j7+
t1qdl+fGC+3NQgepFsNTO2BEjQMDruaYj7JIJPAQPD/7u2VFZeREvzRPme1N91lQ
5e5mFveVN5foLTqCdzemy6dyxX3k+H8ARs4MVm0mvDA62cyUMELnARVwpDgjHi7i
lYXo3NGEnVKEB001J0FQmCPzwkB3en4bm8W4nj87Eti3uhoZcnpY2YiRHCydM3sM
xjtp1oZf0iVYxIsey5tnjqlaoWmmG0gbxj2K49YjFgKC6GaTHrJU/uWtJJDolHyJ
qOIJTwTjhNfxx7UWTaUzrpWRTTaSoI3pAtg8yNZQnY+S+Y9md5GOqg5V3YsYpqmD
Vq1OeOzOoW5SGq34wGTAkeldIX+r9dBzefAHL5aHZ/11270PncAoTtuFlsbGydAK
5iJ2TSdmHpMbVqwdwacmmqdCJFzxvysB1M3QbjTKRmvnSb8HJZ5lZ2zI37AiKez5
2lZju6FUZXXVRqNKir2dC+SpngCIGPZ3hCan968tIx/tKcCKaYSrgjzt2oNcdgwn
wnWj3EwvWXHdE6dfjO7YoJEsk57tuyLmgv+aReLe27x/1GAaOpzhTPMnygqBONVQ
b3OGepTBRZnjnI7eITdmbie5JQa44molq6iSRVmqvogkyjYuQGIElOUPZEXzl4pQ
ETspxsZxEXDTobn91r4y+e5dB6eku9bs6TsCCmD71QE02ANp/K4S2CJO4WdJRmQU
/FDWHhYltvIL2csqx/SBMAoaDUa5z1HDhQTGAVo3B+zFjCaAJjyVJV9JqukqIeQU
WCVfUeoMsE1tf5Ry2bdFhE991PCbrFF/ig5c6AikwnEDT9QzYGRpw4XhjYBlXc3i
nHqgZv83afgoQHZBnzeiBhTRwQcP3jX/f6zc5Hf8+oL1j9L8kKQzeIXd58iMvUpd
30zv3cVpYzwJ+fdzRwuxY2IjoWMnfMAK5RedGdJ2EStn04hdAH5fLI9pjtZK9ToC
ZI+H4R/GciAqF5WBLMhhsW+10lBcP4dfCs/4ylQlClGT50FE9jvFTrwMbKzxB5t7
z4KzY8AjUhSTavKIg6RjaJnKU17V2MEYeAPeZznQY1CmmeULgLz4LN8foD0/ZfUD
A/IIfGat0w9ftDkRtAvheT/1zV2xth6lmLEqHyxYKOMlfG615WKrgAcVkpzI7U3G
QMgToX8irCrMJ8yZzhAGvip2uB2EPiTKVqveNyCzC5P4NZcUyKI9VUxLLnrjhEdZ
YiL4eMZMqwl+FXweB7S+DQKW3FaEC3VEhyChHUIF8NHRMHnaBvo1kBmfv+7CDC3v
SPWExNaJL4/6GByb6SMXoj0a4D6jjjaRJft/wgoSv/urNWi7a/RPb8sqJyW77ioY
MosBJG+rpo8Rb5G8UZWIXQXcywPp4YvDlO2q9uLGI+Dyv6AcbJotRMcd2hNY/pvi
5UDLcgQQ4h9Fi4QLSx0Br/R5uhQaC08XB5v+epmOgWt//gr6/+PsBEfj3WIfCHJY
G9KlUyKS1eolhhiTYelp9c2WNTOIx5qVoVjiD38HdhEMGK9GcVVwQv4FMdpTCo+i
rvqYp6rEg5zOwhi09TTOo7MtOm34LxZ1VWRBbPssLYp443JdGGAVKZ/znlsUtoiy
0GfmZwbrInZL25iT8zGCb5rnJs+0iAxBNes1coeLike++HDzTkQF1sL2EzDFjAO1
IMjZTa/PewO7NO3roQAplU3VCWvDMuplkNims3136aSJLE06IB8i0Me0LHTD0OiE
jCtvzmCOQagpELgGXstp28y0JEJhgiu/6SFFv1TLnRAU9lGr6lSCPDfT51kFY7IL
hhBdjk+lRr6TMDyNMtFuprAwWZ3lDsCfoMiY9iv60gkhl9xPIRMiqYo/Odio0fTI
V80R2SG4HKhi6DfASAjbqfAqqgDFi6I5kFYdAWEA6fYJ7ou4lnFteze+z5x25HTn
72vdXYDYr/uFhWkWjAf+WXKcWe1sPM9E4uek2h0JMqT5/IRRwYXuwl1QAyoZNwvF
Ffcbyop25SkQzrfItNwuoassIOmZ9a7ECeGcV8BldTmOcNf09WCUY6Y2VMp5pZBA
EyqfSt7gKBWa+9vavTMtShFzOrOikkH5dEVWrRvRLJ+dSrxbRcy2MK710Dq/Mffc
1BXcAvJT8MUmWttj8kv0SDJqM7LV1c+6Y09cCnDOwYfSKQx07yPC7VPmguKpPHVu
a9xVJgqcl44tTud5XJwC8aoTCIHmYmOODrS6cGa8btcc2W1VEqcpdYO+B8Q2ryLA
zMoitV/TaevhGKf9KrVpuzPKbQoCUcCMsf5duBtN1I+UlOvLCXsb3lgjXpyYxM+a
qtMQZd2ERyonPhX6QHshRZMzuUDZPB0MuJhed6u94sDPVEYGrs58QXUVgN5P9SYU
Km4UOWLH4TY2qye+SqyQ384GQtz6t3cjZcLkgQgh2cMahSMHggUBYvCj+zF7XIsA
Auj/SqYm1l+tbPEasx0YUgslN8ZFomXOgerT9138e3btfBHUNR8ZxD/fz3R4A7vF
/NyplwgyggzEH0RVSD9RPtQYnzz9Yr+U2wNkLLM235UFTj+pL93oHjjJViVHVM/w
WsamoXtlGoL3Uw7sjCoMLNpiaZWfueFOWAbe4rEhFcZ5AAyHQxgefTOTtNhgn+WQ
nAc1BIJi5AR8sH3NTvyJDCr5i4JDM2V10IyKmFjnu3fYxQ5QedJWyFReC8TkNGFd
fPQeopgTtfFYShX4HhcQ/7y/Vh0cQhmvdleUea8XoTTZWMjuO475/ljYtAxws3fG
6HTixYY53L/zjW2zRN8qW7+CE4e0Y508//UCZuE12ZA6Z2vPPF5ymtUogzZGKaHf
tLk1SLHmHloLxKGMiYg+SuBlHQM1USPBB1++60wXAfVXwt2PaxBDDlePpQygzgBm
pqYBs+hXbpJXWvbnpLlLyBReOsgVPzNpFSMRz7C/U9Kpim+dxmWxKu8Bxspjf1J7
s0vyCuctxrt3kWC1mNWaeiwfz09ACmviWLnF2qXOYHi8lVBrRV52bIWEsfR0aksY
h6DGNOcLwNwJW6zJDkdQAqEMzruBaSrjDpw6708+98aP5sdpQkMxUWSVp5r92SM6
OWYIreblpAaOpqvYGlgH1lgv8KTbO5BG0mTKjcw0Gy2zTAslcfJY0NbP82hPzbtZ
i/CYhWSLpCuAgUzAxUu0osAjPQnSfRKb8JGoFIN4snYJl4Ji7tJ8jXdV1fh0g4ay
DwLX+DNjqVeApjYJ8xaV4cyKf9JXRU1P8HN0Q/gtv+YnJHtDL6rfdrKAlLF1pvB0
d3phv5o+sCSQQSoNahYdo4yRWja8lXtEbZJhhJ3yPf8qIxEFbv5A+NRvFiZzny1M
3uGxmjWQJWockMgOaPiHqh9mbqrO6IlhcVMrhvHv/K07ZmtuymrkG/u0fz7C7O0Q
JcmK+1+Z6CWn6SYjGJpMZrj++NuwB1dQ4bSsOMDQaioQ2vgrMxXvCjSXVwMfdEpJ
ORAaw5Vuyi2p13zNO2LIjXmRY8KvL65pjHF8lnJGjJm9eAsfZa0Dp2hmNrdsfKL3
sjagy3pZrpGp9p4BL35mFnsXG9zg16WDc/GXwEOgUQUvur/XukLOeFXAhs7OptaX
PLVWgijllFZvrBdxfRrKydH648PWpuqizx0grEFGDW99Cloi/1R3FiPD5dfE5ava
0mc52ABMEP1g8Uf+yzIrk3o6eybD8DN2BBW4MyNfT8PtXUQ3MPZS1YAkoqy6KYyR
7R6KJgrmw5EU6Eqp9r5s05PGRS4Fxd/PoUy0e9bz+TjjcguDTMA9zONsmzz5poQs
gqlTnhCmfwEPGz89Wp0WSa4c/6WAfZbNN8DmC0AYXWQNQjRupqyRl8wYNcbS3PCh
BYdX+5gWoTq8IIM1fLKkBw1EiqwB4xxVhyJnJkYZ/G97p8C9H8dso4jKoJ+rEXM4
KyNiyN4/N3KZ0H4AR9zscQ4BUy1jq/btOqr2yXAM0M8cWRcFvLLTYu9LwtNvbDMc
LCy8sEff6tU9wTclcpkWcIzLcf6v4USdjUYOD0/Uy7C5ZRblAnS5r8nMkPNzCqW5
ldsEzZVpjNKb1zQEyYxG9ahI2yK4TBsMhAoJJ+OPQDt06BFHSDbYwptnhm+gcaB0
QcjPqa4O0M8IxXc8zD56NO4yIpV+rHqcXzIQe0K8PzD59s3RulAdqznw/0jjuqrg
wMJqxKY1U2dmfcWVtnMhyroXRklq8hHxpRPbVhvIoSgA7mq27Mp0szdTeqpOXdJA
O65sa1Seg8j1Chm1rTFCvzwqMpcDAER/ibpbPaj4dtiOI7TJSkK/0+v/gyUvEoN+
tZjjsDaJXhbYZNfRX20YoUPSEdprGX+5sjN6pYKNPH73AWyAWvsfvM+3+gNYtCCs
Jl/sSEaiB3JHjuvo5WjE+j/iZ77xZ4X2IswaxC1yWSfSBSPX2lOuyCXrlqhM7xFH
xos+uHoWbzO5aIpRbWHGNxtrUvGTSnnwqrG3n2uEZJljN/5/3JmnoMJo9m1ZDXbb
XkprTyhn3rSA14Lj11e14gisNbbCGZ5S20fLEB1zvZl5TSpw2eTomLp4Bno6pEXN
5gE2hfuf6oP2POhSA8L/5qhtHsl+uOWQ4x11euboQYOuppL3ZEZ4uvCrz3fuMylw
RhpH4AxWN+gpDQmCZW4OCoRpCA7IBzeNm8CZWGQKKUYROQOv03xpANRQBsvnx3X2
+zlegB+tc3tGw02oKO/ZXzXxDRD21c1Id+W/+0Qcgn0oXv99skJF1gpidGT5YfNJ
HdIYcEq/hOU1mp95tgfAlBN4s2wnH2d3Pvd/jpr+lO40lS3ZfVF/rnsjSuGHGQ5v
ETLdfFP9chNr8ao8dyGlKbvaFVqt/4f/Tq8OH50jvzT9UJrsnnbX0VkLKQoK+Ouo
N9S2K7iPMOyRSNB5kyzfTK7OtkZMpMeQWRn+/w29rzmYk8DF15tzEJ0PjXP4jRGt
nOegasEKVDQ8sqZ0V0PD160uKBKiKFXOnfbBcobfNpIXNYcGVmJIGpkRUTE92Z7K
dWnKHXvcFnNtFrk0NrrRkcILodfWxTWletG2WxnBuLe7Ud3EyZGhDUUw2+eKIjqq
VXYLHtWJ+4V4D47qxj5hQpUQdQRlcHVeN1kDNWY132xB95B/RZUXwh5wb+Fk4/mn
CP1ZkRw9LkoHNWmUk+4seQrDJlADmzyGwxaYTn4YJ53JYZvDqIxFrDJxJMkmmpp2
Pjynwv91/TmQCxYy+wj04DFrLdfhwhva6ZxxYNeMpsh6zaiQNg/8zY1dP0CL4DmO
xc4ioxqiGb1lbT+vXg5XF6gGOotCPdldSFe82/JTvXvmBEpUO/zs1hiHBiYyydWi
pvh+pZtUzoYADo2llljIfCF5HaiIXIajhOR0JS26hYsU7aV7lly+MGyuaSaLy9hT
OipUHlI2ktQgTNkXeZ+znTfydBkV/shYqIPvsSv7s7U93yLBKuDSc0BTJkgVPdaS
kI+Xkvu83SeIfiBVNwNhzwSqAdNakCJ4ugmfdyM91qv71D3VTxHFbayyrMPiA7bO
cAMQ5G7ej8IWjbMXM2diy9lBBXhlBeGUpDI9eVjuT7w+B6GXd+RUitOlN2/Z2mMN
c006/0DrqhUuYf4WqvQ3KTw5b88rtk/blPDcxToavTrnrfkbMHPuPGu3Pz2VFTT7
BcDO629lZvlXIoagpx6s552Om5FEHfCTUuKLZ145tUlcgvbKS1QI+ErFs0zgud3F
a2416S42H/nATKbYy+prYg8FWF1EsLJzmI6eb9/snV0PWnIJckz6rvqKUC5QO65D
95e7fm1dibapWbzGY7xWyornJsp4KzyK8gBRgQjs0Fr0aPRp4zZ1rB2DLr/V4koH
wCZmIEfFcC2NYWumQRmL4mCa25JskaJmYBqnjvbNOh/QNW7/bCkbqsRyYROw40sH
p9NTa4KNrV+e8rpCbNwl2EQePFo5n2TYxkNQw0loFreWNGXF1TaWwL3H43MYWV7/
kpA7cOi5u9SzfGiFLDjmrfg7xoBzUlLkGmRZEnq+Nw4XUy9U+VOCAfoUOfxULyug
dAHDTSVX0nh12Ie1lu0PWJlMbo6MnNJ5tkyYmoJSiTNOr0rSOYf27LKJNJ9pPRN/
uKB67AaNalDU/Z/YKGOAEN61z5e87lCl5ucNjqJ9JXLeUEJ3+Mq+sdOvPMWNwTc/
nRZM1m6l83vCd+sF+c0sKuHL92xt3fEN0zVL2mVmiAKvg1sEEJfBvAAcOCPuhqrt
7CzfAPhwbKynmkBeKiP8Hw4xtBrGXh4lGUof6Q4isuBHYqRPbAE4ORsNE/eDG+M1
Rl6T0lktnyReddrKCeC2ZzXW4OCvjiEBBv/JyDidQmtObDrv4yd9d89YCQZEk8hR
laGu5jI+Ao5NZF7yfqbTYfAOjLkl8UpJwvy+MwqfUp/UjLxLpcE0yJgBshjHj3xI
23LG8O8XHqN5QGN/75XkYNDi2v+fILlmZ6EFHr7ukRrqCR8hQxd01Gc1VqpRV7aE
IkTSf7TqrniixvyF/58gjoOkrzRK7txhZX3VGq6SACPAOgc5w8j7IyvLM7hiqv6s
YwZO/f3jTAPL5o2aIC8jATMIXd+IH0XVGRxYVvsj3+Wipbmg4Jjsb+rZMQz8g+au
X4N/RY8SGh7DduUgcjHEKA3iYWKqSbSFQE7/yMkprH10KRRLfNf7km4yJI0F5dtv
DL/vtGSrZ7uz5Gz7b809290hgGhO2iRgx7KL2ENf1ehPQ2k6VhaCXi9lN3H3zsvb
8T+Cl/QWvuF7xIR1t5MYGsSB9WeSh3+TNSlC/jkQWlybGfnIvl2dbqp4X14J7PBK
klNlM5kOOt3l+KCLi5xM4qVJIYphZDvIBJEco6Q1P5ur/FD7vwAqhkcgun0tg/Bx
dCKEXUs5tJhoXvRtJQ0v4p7lcjxGD1lOJtOHD1gcktKMYdhptSsurygxTohrQ0UE
ZLEcv724fryPOrOcXZ/DwDwfw3mal9yST5E5QTah8+EqDXVxZl/qa447udXQEjmG
noP8kmnKghpK4zJwNfM9deeQEBDfQZ5blWqGEvldOc8kPBwdmLddENS/ucQek2uO
iCCFpjiFEUKqGp570acvk+yNDY0isvbpQgWy+4/yt8bG+pD3Kx1JX84bmyIrN5TJ
Q1X7ZjHWOchDqmhQQPF479T4akwkEThQtjOV+/0TyTfoORMnuJpmu+7fDNW5WsVB
d19m14pwGQfulkkT4AlEgZNIMTXgOBHSLCdxR8GHn3/zAmEftGO6S4ew8pvVOzXY
sMEQTuLvcAjqRQLEAmItrnW5w3Ye6foGYrxDtQCe45MWpFMeum8mehi1N553nbNG
ypCIzq1ypAyOA/1PyhXWCMA0ilMfRgC7LCATpF8ygs8+wc0mu68PRYiqx5KEpQfx
pBb8Mcfw2HCYVLe/53J+bzUEFrC3AFK3bmPvQUQXx8runa4eO2mvuUUsfJB045Eg
l25/G3ySl3MW4o3/JIK0hwJI//8Go1BeYgyGxWensu809oSV/E6DwJWSS+kbJITs
JIwuGQ/thSfU3RTdSiSCerncqA1zSLb6mJubHa39vAL0/3rrxxaEkhf20oCAmuNF
HfLLqEidvwl+6UbWKuVMsQ3YNTdooBMNFl+BgCPGeCI3Zp/IbgwmIAhmmIEIEnEX
hW9qjj9TbOCehL00RGKXCiLGMAyDHrVTrF2S1dsWU83/CFPX1QusL6koJ/Xs4j/e
ddXHrWdnapVEvpiNiEm0XZ2jSf21kI3lX9z8f/2loGUOXSkjSNO3JcTMW1w8UgDL
N15AHJngyYSmsI1/STc7QW+xwU1/utgHSl76oldXnbeJYe5QTCIf3jLnGt9qFFTf
sUSXW3g0Xg2fKsCATaGSig2OnCMcmwYCevmrRP+cy/tPacAaNwmFnYs+m+ozR+pT
xUPjDSBpANrzgr1rkKrbw8UuJOVUyPFu0ePiJHr0IyWufmaZB8FrYGByIJrKlprW
PPcPGfAHIn4j4LslFAASBmjFWaOhEAPu86359tVgrwamSG8cMM7Q4rwsmcNu1hLT
E/NGLYNHaHiqomYD/db7D+QpDY7rXfr3imi+owRoLE63BmSWfQG+5HLji+QUyDyJ
ffQNfTCsQUab0s/Om9rrbq1TnGGLyt82oEpWr7mt9lGtlHfFYZ71prvB+I22CB5U
Woq6ApWVW5WiI6bt7VjyZk+7JA9YRxgH2O3Pqjfbzk8nUFBwNfZNUejYC7+Wcm20
ZC4tGX1hy2x0lz7G35dqyYf+rmV03Xm6cWkP+7dbbsx+eSRMGZDvNKXZ4Nno55eB
4yLLNBAGmUkbqJ3RTiKgEq61HbGZYz9EpUMG3/IMLZOmXQb8hWOdiERJseiuxRgw
Kv5S3tRSoTF3Lh3cm7SL+PNIHmvFoA9iSqk2lbubG8YdYj4DpafAwNnAu1dHQY3z
Qnn9EbjH1Sy2gRUz3qH8IocSSn03Rg35Reurob0Nl941T7owet4MHIVaVhmWD5Iv
gmW27m23Z73+L+NgIb7/R2j6TMbANsGnFMLPSL8e+005F6vNXqKN2Xpi+oZ+pdos
I4PmUNhqJ94uMpFIL84Rwikf7MbAPSqge+QQN20Drfpumo9O9hZgU3Q9s5nuCv0W
3etYggeugUNu8K62ozIVbVWDHYy+mk9XlcKiNCVtMx3lI5nUB7Me50uiDA2WleeC
aim4KflWGxXoBqzlHdBJTP1aSp5XdNOXvO13QpciJxYtTqWBHEYHmYyxJJdotvyN
n9KdrUdbVOLTMg+XsJAfLNjstT0SDBiyXY3/++yWLH8YdB4lAxbM/60L2kgsieZ2
OvWjPgtekhW85Z8qKDVmRzzJBAhpET7TWiXspAzZ72hWWtlCUjNcyaoLMYg7pbwZ
KmomS5qara26aKBxJ0KGWHFD+ZJke4TRcKACWbTPdlxldRUq404g2FK6cVIczwKh
amWMZRUXfcx1hUUloF217pN/ecsjp94QCFOO7jGAPUxVDfWJfsaX3ERQxebrSZlV
JZFwd8Jr9ivzf5UgIcclkXoSGbRpwZ3jaBB+DnGzqrNDuaTQBKA3Ju1h3hTYBz9C
EcOAgy1gJ7i/4OhWpdaEfXXoi52n1jA0c29KSAVV48CczEbh8fQbYJZcuVYyH3D7
QJCBnM3CTVlUez3lEovv8MQ+x/X3lFTJV05LdX/dfKmrJNnyebfC+Vrq1UpkyaOA
NYr6nvmaiIMb1yEDnwWrrheHEKRZSZ/umvrlcsgemM0saZhgfn9cWPozeIBqNwuX
3rUpeAwSnEvJubcC2O/1HYXy04Q8FFtFYUNoN6udXiNXGsf6CckT4WMIgRqoKC03
GlN4e7l9m+AlsxD7d2na/z+bvLi5tdK8hR9yezo1JaKGR7rhnKS1aKt/xR9vt7nS
XscAZ9UoZmXOrrUMHAkka+Sjs0fRsta+9hHNojIFbMXllA4uAgPBhjtKqjat5IID
+88E9hbkoOuAUSmyiAEL1GmaHdNHgYSSs2naWmXpKSG1ZODcJ4ZWp0Irl8IrieRv
EicETOTS9T7vzu25Bxkmo4gMvmksusnbD610YfWPR/Mo1bv8d576MFbrfs80tclb
FuJvx87ZLeybJxGjcHhIxRKsEJvR2SpmdnGLKjg2nkReKQVJ4KWzw/3cxNwAWZ9l
a8BrbFlmFuQu7vyw0TQffe+NHNbsMkt/h5a9id67OWVevGpEITZHXegKKijK+S/3
uVFzWVx16wHPOjjVtHuTih2XG6Ut8mqNrLQ9I/KBwSM7+3KBfOE3wPIvIA5T+JI2
Pi60Q5TSFManZV0m2wwUgE5OAarNylqORerdW7gnY7pxMnqTxlJ2UYU863ICJPhR
RCNBiBC4kamlfzZC+294WYJ1vw0LquWutr38hrjbaIkBsOcqUk+vIAZyXp0h5ARz
h1dZNCdsDpl19LCm6IfP7BMM6bR9H2H+iMFYWSaOtMzd4dcM1zmhCr1NZNlt09eW
mPabVlpBGfsUMQqiMhdfp4lgz7OJCju5OxREYhDzGR4pVOViZPfcsn5YgM9BHSW9
5NTWuksLjH0GVJbaNuCl5lvYgKPY/xv71f5rF9Tqh2WgPnlc/xqUR2mCcSAO5gN8
V45wn19urWOWqCFhUBAXzOBhBIA2cgF9qBcfbWKdQtlTHKbm9rVZVspAtLj+NCCp
Co8h+HAz1CLN01Kk0jhl2gcOBSzf1i5ux04d7PYvOdC5cG8k/yknQlLKz1zFT9Ma
zdFFG8mMFDyuvIOCskz/GqrOeqJO0TryIa0hi4/YFZnVuWR78RVrgCaV0VCdCJtZ
btNTrzIq0sBgxLqqH2SZb8Nauh575Xq1O/xjii0GdumnUfla3u6D4aCdfLWn37YJ
WIFgRIEGqlJutn7OP31fT1yIGG13we0A5xuMoEZqr9yz6zMVwI0nE9aTbMM2ZhCT
LI9D9bzeWg8v54FHwUf88xf7VQnp7y+isw7hxwYzxAlGUtfaNozCy3J97P7nhdue
Au4zlLIFsthk6e67rMauWCKCvWwVErqN1obfv0ZKHquENgPmwJqJ6OgVCMvCsdFY
EHUono/xDSVJb9tdOD0dzt9bD8Lm2ss4XFeY9CO9787K0bJQYpZSctKb1IMr3jZo
FQHHHFOwP+gxa/oDMQccva0TlCyYxIJBPQZxe8wKZVmuQF7UrZBHzFeL8smx1TEI
VX4irYhM6FdWEH7y+mQqiWm6q8iKvT0NE5+m7PKKX6+fPvMb69sQEax9htmkMGrI
RCtUlL+24XfagSSEHY4rr/nPo3C1giX7cmPWpzFhII1yrE59ft5HTfxFR6w9sbhN
zayR6IKhqMuNq2LxwzrGBa4MrqPPzELyI8wh9IqZ2bWYxLTU1n4wLsv2wSlqPuga
EVUboo7cU2JXr5Ukut6+y1T/zr+5P+p6b/bpPNhwrU0YM+83B8EVrIcERv9AYX5K
sBcQirrqLBQ3GuuUYZEIHdyv6r3lw8Q5+CvmYtVUkKFefpeTv0bpxi8xBzCm56Ab
djNE7WpFDcYrs6pvHGhUMAYzSXYpXwufPFypgwOSad9bpBnqy/JbQo1CxEb8g5zz
dpO7+LOlnxwEle8bZkME/W5eo6M1ybYoEd9YaMJPvb3+6mOZzRIOpPVFDQhnMXEB
y8pW8qvvnzGO/4QAIMA4bPvf/+JIvi+00OQ6lSCFxazZSkblUkr+d+8ToRCtIKKW
pe3XPDnMl8Hs7F0DnTi0aKEYPAwIb9LYspW45iAtwYpVAWh9cU2f5dl5uP+BUxFh
enkqfXuHGUFv6DJR4ItUFd94t01HKfDFlJbxJ2KHIJSOn3AYfLUl8bG5c9Vd5EBt
VzyZVkDsiFVWSWbEFDBIOwjsoS3O0qIo7dZd7zY+ipeYt3HGPkPA3+/53l1gkXh7
YrDs9HQTvo8F7GsePsJKHHitsqC6I3ZGH1B4ik1aGmD7ICn3yJnLb4LxwDIl1Na0
2Gl79lO7TkntIWaBYvXeCGEO7GxksJFhNWm/23Bb0My88BxN03ZPB/JpxINrS4LB
XROis8XTFzJ31KT7KvPicRnre0Cmn5wZMqysI3b1VOiljU8+vy3uZ1R2GFWCQidZ
00tZI/AswMBnfQXbBNkHLapYR8OBADs5RcfCvOxJmVRiaksyaeRcSbtqsRVIOky/
OrMjA19ApHV0p3TCQwTjM1P/WDvts3ui+QTw1NpELbMvRRiqVPAS8Kkd6oh4N94A
QY84X1DPfhTalllhNw8gqpZ7MKvj64XtG2Gt3jL6XqwgIR/k/UwmF28BQi2fej29
/Q9TArAyyO2o2wHsgDBuM8ZGZxtt44YUs2PIVL0EGE8cg1debMCYXoCd1P0RNLVz
2wTcOxnrPmj7W5Qz5c8PVLk4NPcq2cjaPjvBToQvUe0wvwjHTaw5fMMIoCUEzfvX
cB3a2bzU+ZtX6cVGaKKXlQgjLYqHLzUIu/P7Zutw7OMLNF2oy1Xg45aa9wt77Qa6
SHgBqfca2d+YJW9NOJ/UanGIAJQP3lw/KmGJoJWa+CxnwSMz9RAV8eHBfZXM7UKk
i3m/isakkkCepx2MjaVBj4mtK89DSTHZZDwPPGMNdLb8g6GBRSfCO82fqG9SY+Lt
0Y6BDabWxfcsZZXTzHIz+gGaFYVoDWyOJbuBl3rieZWt3rNFmSDGJSxMTebnrBsB
MXEPepaXHU0F9pjcVCeGXG9k705kLuniYrkrVhbtSIh4E7JhMawP8ZGDOsYzEB+u
O0G5F0yR9+TQWuJnug37p8TWigQsdf9yl/A6duQIt9GxOO2T6jqKLFrTeEbHujSF
k8V3uryepj0UP0qsOv/W3hFTYdOa7Br+6d+DWl4Es5+Pb8CSlTA6tUyLbwiUovtL
Dop35AU/9RnLTND66IhYY0HA7fVL9+xIkufoZDPcWrcQGZc0US6f1swXFAHeOLtr
MxOu9KJXFsN0bNyQzkum5U0equQBU2hmwstXzVuO3j+Bke3qz0mEKS+D8F9DcTeR
HqHOoX3Y2S0KKBNmV1XCny7XYndvl7WuNMuwTiBZ5wgLe2sDN+VQQZGnt2NA5EoU
CRxrtpTwpxULJy4nnEivoGXYPEwPxSbGQRm6bTSrr0KukI7ZO05rFOOo0CaTNzWs
4EdCBClQJ6hgfS2+HsX3JWHfB14CZz6u2PXTsYZZQixToCAI4QEteiPkgmyUZBTe
+A0qrb5fmixlpfcMXBWDF6TmsUqWGixVN+BiK3oD4XE3ZwMjUSbjyxF7lFGq3W+E
drHOkg9t82REJrMhj0cNSCLkh57FsrlsJ2JYQzMZD7ym/BE7ev/bHLZ/LVQUh7wb
7PKXQzgLRXF82QlHcPksW+OAN9i8HWCWNn5Uy5I/DOktw3Iu8Ktp9yQ4yf8munbK
OsMw3FnkdGnlaQImxAx/jAGjxVfwzy30m4Bt7Ylbxfaa/alfjJO/YcpPI3WSXjbv
LWWRLw+8Hj3nwRbeSk7bQ2nOZitLbg+4dTHSyRAq982iRI3hMjAcFoi5vVUo5+fc
61PVwbbPherWOTTyZS4YoR+xa4NZ6RkI9uABiRnJZZRWktXuh4HL8uV3fBvLuLiD
l1A886cmJzcikULtecxQ+f7CbMLbEKua5LtJf9uuPD+Y+iVAXxJEPsOSF1stHbRd
3UK3EJqUwypf3i3akqWTp6iOc6Mk63ILYg0hK4iurtGyNTxMOW2j8bSgvOlYQTgz
/UYeTeGxljYy2HjkuhTc2C7ZzuHHRajbnVd+vJpJRuskSxyz1rhyPvAqc67/r9sV
63oiP1Jcet/5MujK+hqg+vHKaagE7OZ1QkvWlhpRZ48Y56LPnZ34fuLI3j/hMZ8w
6At9iuBUUS76EISIEkuMPvdsCc4JRcan4on+7qDaFyafFTwivB2qC+GcZ4CXmCrG
6uROp09ebmnpxAY1X5f2q8YerQR87utMGFLKq2SA8zN46e4J4fi1I9epzHz34Zct
d0om00UR/1BIiyBKSzGhLSh6KTyi8FBE3xKN9Q1JBIOqnfYNxxI1nBZeuVrH8KK/
KJ0vPxWrssC+ZDzMD4EeZW1WEukf6ul0Stw9qNJVVHB80t/7ga2Y4qfCupnC/lb4
W9sOCXHYNyTLG9/wqLxpJX6GKEYUegdEsdqQfivfRGS2imVgs/2TamMzyIvRZwPT
HwuMGr8lUoi3O9HYNDkzMRlNqyLgkmdSu5m8SrgIJH7UKKjT2eoCsXCwO/i2EX+B
nC3vv1wMjzOna3Zbs5/Rl4FjuVmrsbReEYV6HioIxhYXe0vABqxUSi9B3Av3sDgG
0LctctKph1ajNCyOSNA8iR/jP+E+cEjx4laBD/LUgtu1r29qqwWNcr5GM8o3pVlx
pjtgQJKhSXZRuhkELtlAVqfUkFcSZW4Y2SIQWRuOrLA1DN8MEbMaQQlWLYBXAF94
HhGmx/Zx/WPXcf3O6ncCexi4vVp2yvmeDLafVzwtyvDzfiswCrXFIlU7xUJu5sAL
2D3QKqSbJD0ZLT2JYfO9cYxrEGerlS4d7aMCOA57/SiA9nVuHDgD5oL4o6MwDXU6
a7PKGyCfOxh2jQTnKD72dct+wBLSovjKF2zKfLnSq6M6lb7MtqjMF0l8efEBt987
uVdWVS0D+0VYHgc58xdYnhI+rwy2lCeURCgWe7BIh+WpE3RT22982hb+bJ1KnK0H
+IoJSmFN+bQnMcG4Sf70kwEFTWPdm4YmEsMWHuVC9Cm2NxzkLt4gjqV5SSxPzpmU
QUwIShTG+0EQ/B5gcWfwsBWwwWCIO5vlstf5eCcMxV6kwyicO1XNbX7FWekwUn76
inG4UYnB8ZNSA+B0iJCY9bpFfTgFxHQdx8bczTV7yoLC18hpZX8X8Ey/lDJQmmhC
qatGMk+pskJftKrA6hvwsUeZxo0c8KVri1CWRvnOpCMr46Sb/YtGcn2XTtZ9kZ1B
2VeiYM8APefy7TSWHFWbY3TAtcxmIHN18YqPzxojKgU+tMBOHWfu3Q3qhBVVmM8k
TdMhDR1tFuewi8qslLYUXS+xTeA2xD2XhPYSPs2bTsxKceX4fNfFbT4Eo4vbhVEQ
Xy2VYHdkmhCpNQEgIwBaOXmoguxFu14MgpbD4xpHE6vOj2D0oePoMKgBNru1Ng8p
4yYHyfcgEu64yJ0EHdtsPqVxGwYbzpUQF+WZ4Ss1fBYKjAqDRszfQ3x50fgmCyKA
3SWlZrxRZFau6oGkqmHThNNWDEaeIRtLxY/MT8x/FsWgvLJ8BlFR6BU7qwz4WwnS
YY0uFyajjsMe4GTYH8I+WB9MluN14mvv9okExQxB+WyK46/BzABVyO8SOIeqxiLT
wWUH3XjM4/IuGViKQyt1C5uD6M+5XGK6SKb2fgbP+3qXIv5EcdT+VYCuAQe3iBgx
fgJXKONXBvvyIfNbtzGF4JyReUWyI7T90iVWiKgAkt8EsMfRl6dQ+iymyriggKFM
NpXFvLJP9b6psuyLsuGWOIR5fwi24lcvSbcuI9wWwM2DUzc9b5AjQZoFTf1k8JJW
xEfwK2TDxUdB4wmu9D9PL/NxRQVcLzpg0hd41y/kLy3Dko0QKUBMexpJ91OsEg6k
ZhBh3Wm7LYtNptUjy+hp5gSEaHri43fq7IP+9YOgDyOexz/mNcfjpLpHCg/VJWNK
pdw/NOVvLPy36I6t3Bun6oh64lT9b3g8HEBaT2CD2i7t1y2u5QVwiDTtfujgD/TB
6d14FZzX296LKkwlwlVQL78QSvpFW1wWEeZhvMG8uFRjf+1JxVJHpSex9L8w4ljZ
bOgg7Prac2dqpQIJ/HHyMtoiLSGtoLjW8Me2GGK+GRzT/XwdlHeY2ZbhV0chUNJE
vOPydmY79JUB83BOxrAT17jFDbcWyUhLKxXh5SdjWGJ5A3Wb8sWE6RyeKzcnbPzV
v5PIzXjNhDfluJh9MqvNBB5ye/xwX1EHzrnV2xTdRV/tYZ53f4e25egBPW8tvAa3
bJ7yxb7VeYsdYwkSuE4iengFV5BUKz6mXT9DnWwGZtBEPo4zijO57ceqxj6+n6Nk
t38PsyrmbFkzzCdk2AzCTaBqch3wpkA5Lul7YA92Hqx7vOw9UvIvjx0nbXfMV7Qm
12jUhCHmDGzEFCEe20Nm1MDX27tP/xUrCn8ID0oTMthd1sFXz4BoB14N7HStymsh
3eGU/pzbFDO3gzd0Ew1D7jxcHvIobkVwZocw68jEVlcyiCXaiNHBL6b3CRGbtsPv
ssk5QM1I0mUf7m/0LBA8Fgk/RTdHX47uVCKD/T2AyhxEMzt5wX+TIL1MroOozaax
HOki+kI7+uI6NZskiRx+xoOb2ImN9v4F95On9OoY3K2+gbg2UvOwv93WW2ryBC2E
ptlVsDvGBPv6qkPYW0N5+T6nnIwhRJMWw88x+HEg0qEfAwIpk92Ar6ILJQ0p7yBF
rRLst7kZ454wACJNIi4gpP2HFrXt6CPIbafD+HJAU03zqXux8uflAd+OFLXHwtf/
78CYHWyQzY9mqGeawpq4+cXAg4kB6xb2DZoRsD/GcHoYXQtgJ0WuvD2PKF7Lsejd
wTCT5qzH/G4tR3Z2bWEtTBvDraIqz+EtMNbdDWFi/5BBB3teWdZxVZvXhVzcevSi
tsQV9UvyNp86+kY3R8NIVDCA1Xwp0yZYyHZbhiiCnT0LDH7Y4XrzX+LwgPNEctiC
RSd8e83+m+I58sRZ2EmPl/Sx5YUOL8dvNJtHxklVcvjq+v4P/TrDrMg+QRzkXvIS
3KWKjdarE9gbpV/i6vsH3p33sf3475LiGq/uzUCjiixAQgIqRQ7kFbvDoU3P3XQP
bglPUD8cBM78HteoZPIvxQxMWfcZBdIJm01Rt4orKGuCBz8ytWVE1V7yQ2633H/k
WOEByfV7Adn0NzSuKUGjY0F/FesWNLLFpXRj6tAUTbf/VA8D5SIz1S/MK2cqLv83
Joso0+cIfyw0gsvRZwa6JgkGrghu4A6OUZPBUr6VgL7orAsAFpKvXofNrWVNxHNT
/OZNCpTFRDdtiFuBjuBfd7Qe4oGmpbgMTc54Q5dYK9CXSC6jRZLdd1XC7LmbDMK+
aD1l8924qF0Pf3A3J/2If0/ELrXw7Box9jmPBkqXYa2CMj5YhhOJPNRYAi/4Kyl8
qN4mAh5Yj3h6n1pR/tGQ2bTKLG4+hP4Zoo1oi0dUTYHxZrkk8eSv5REk77NXCfME
Cpm30EaTlF8WedJP/usbfypZj7I9VPpGKP0i7V/olGd8NCtTt0vl2Ww9IjIMjcUW
TuYYU/myECB5r6UPnUKFhXBAOjyjlwMbs75mvJ7thuP1LSBwzQ1SAqJA95P2B9C5
rryIKdg482MOu5HBPDBKIoWmL8znUSgLlBfDMWLJB07vFOVvNKeOCxXCSbUTmwt5
ekVXfWGNBpD21Eb8tqFVTDTRfIuDW4428hAz1smrFhZIcxlaC2tNZELYQuwTqLU5
EwJ67+EXUw1zt+B1RO5GsGDBDR+m5fhfqojIU6Tn2QoI3m1q6DNNAukSIuGooaXk
tgK5Ktzy+xEWxlmf/k/vDwKyau94leqBLyGkyThLsT7pp/l7vBAzLP7ZYDQlabxu
HtGFNdHNx8IImrl7dJ+7INO5vGBqMIj5PLI6b0bMD92PX/zniT2DMVpAqC5iZ1Up
QvDRTiF2D26atv2i5x4rH17WXojvSSgo9mVtO9bvSm6CtuUbmXkI0ybizzWvHhpx
OmWdFBKz2ZbzYdFQ3ygm6m4Pu1wT6h7MsMYH587w2Sdy4MC1TKlibcuD84PgGXHy
fhmJ0aHI/TNcj5tXC6vfsprAgfoh9UCLUSW2BdJ2U9fBEuuTriMSQ9vJswb0tvBT
ZEgSVKtMmHq84KJXg2ugy9Hh3+apl1Py7IC5GpACtP8y9oS+kVhqJ+8dMZcxtATX
wb5ywVcOjTAPEzhmR4PLKNZXkakV4eskD5wgN1e90+4DNVJ9dHC23p+2OVjCRgYa
km+/F68dxKONvlPWiGutGP+E9ewDxFXjfyHvODc4JCThdK+CqxGEOzXStaY2ftIN
LZN8c7AQ3uQ5uPfmh0bY2TyEvS9kyo7GMQBaOi5syqfdt9E9dQhUhs/jmaHXVG9p
m+kijgTsMzxbO0kOhFs8Lmaczk4S1Bz+jDns65xONP9oet7O52mGOvankxrOE2pH
SKZdVJDm/27aRtiqBTnad/u+C1w0FMGbZhaEhwO43713LvgSXOudYBclfSegEwIL
/Hf0zk/wGoTu2slT8a4KbdCa+NXQgGhbdUdrwZVnPUZWBil/wClHwR+QjhH/yWn1
PkNLTv3ae91tGee0Nt28V6Kp+6r01BLVIoOeXzPiPatdVs7s42OCBHG11PJpiix4
8/94hRFuKjUitZWt9wBZFsc9S0UIFUeCZetij8qFok/kh2mreT0er6TBoonTNLr8
1PXhgVvTkFnneHSFRHVo0GX6iUApY6XKXm9dxdDYd9fs0ogJTVaS7/J+i0WjLp9b
jTu5pGOOG+6eA15/PLH77d5K1EPmsK02k43XMIbgc3SJ4cExodLg3be+OUj9172t
xtXunrqLFOqMAOzMHf/xTax/KNke5vyNDogndvf8Bb1O9HiYzKmblQ72cFt9UoMf
5DHWcU1MEy8+rXmTJvhTuFxrHa0LgKk0oLT53ZkUCk5sETZKtbbqbH/+xXc7MgYT
lh4MONn4JTmsRlJEYw624AqaqcQWY2RyHaqGi6tp1+lhjei/OS4mwvMFvoiOoDqO
NFsTBBqHW64zAttk1CcwnjbtgyeDbzCqsxxSYmJ+4+zgNr63E49xzfuavvDzgEnJ
XBblifnKPrJbBeOeWsllsbZHCUW+BYdDFTe0OFBMi47Gp4UwOU3Jx1FFKsN0EYbi
tIDH5hoTtgF8MGq/13qWexwj38Rwzjh478/tl4Oyut1tgbn6WjNjPYWJ6cMxFv5V
vJJIKbvqCI326oGZiblH/P/7CHOdFkhdkAkf5VJcxeO8AWXqw/wSVfDgWijBa/RU
2i0559r+5Ek+qjkvrQFfzJdFp7Z/LLAltokr1a3hBzmCRsN/E69zL85/x90PYAGZ
9lLX9McQLfmHqDJjDE2Irgvg0Po6SMfr+LHuOk9l/B0IvsHRQeLQapiF2TnRyDsM
pdd3Fly0pPY5nLU4V/z6/s3pYxSVFjx5sEj1hpypOv37P9X+SH+IxIzYCT0vWwYo
TeSTZwkCAb5x3aOXr2AlnrQzdOltzVlDtv5PCGtsI1M3eoPCFCuedeb+TLt22Esh
hOElsQu8tWTTg149tPauYUoW1JZcg3Ay6tFsY6UvFd0NYlviFebqqF+3aa8bzxJE
FLLlCL0tog49wrZrnE3G4qNeMlNV/ilg9diMnA24aNflZ7zJqZGB7RvzMFiCV53z
YdSATGs2Tg6m2JNn+vbbCRte3ZgJH8OKyXik0Vxt+3k+T8I4Amtrngg71OACG2Ab
HClkvFWEQlPSWp6araXnh+09PheVMhF2zAUfH57s9CE1eu1EcA9YTRyP1Qc7uh3B
9YSZxyGL3iVnAt66TTEHw/9Qa8pSTCOCYCWdb7sx6xyDfrEb++jGOcAIltqKetrd
1hTa2psSZzz2SuvHCkvS97TYCg1/B8dRl8G/AellCbu9lFLMcW9siy3Fric4wVIb
iM3VOHHBGC5hjOwfNs41+T/pj6mbf/EyeG60o3cTMNfh5ppyjCEi+MHd9+xLyWpP
U406fgTodIKmIAHce6L2dxg7lwdGGRAl0H4iPt2azQS+EMRCHzUByavq6CibCobu
GSv1KQOQdzEztZuqjmL/4bFPhKHI0wxTZiJgn2bFyRycrrpp8OhwzCsRwmVvzRf9
IMXAABvDwiDnCTXSSrMkOXdbKA0jpibyknzsBVkT2wTxYctAKxrlCPGm9L3fR68j
6+c6293YCBiWo59K+BiSfMoNUFGfsQMW6w2lpRIckvSxFB9iiXcx5v8AE6N1sHNw
5OSIu+s0Worq6Vwnwxq735wmkaoieliJ5g6lEuLBNWlqkWuskdkZpK7Lq2bhNMzH
QIcy4EbQX2bZhwh41AWX6ezGc8YBZ6kgpq/T0a3kPiVn0jEpe7x2isQc2RMnu4l6
nrVhJOswhY1C0pWevTnIECbYZzbyoFu/zdhkGeWCMUnD6z9w0N+e2GWFfaVc0wX2
4BGRzkUpfmk7Ef+aUDKyFcLthIGSxIKzkWfIEvJ5UnreYREaw0ef2PoBK/Qf4f9p
8ahvCdh9mpLGk2IwbYPeVf1LdGr+iwSgf2rvtG2g+EUgmBNaeTSkjjNb8OKt0EV+
j6GcSrw0ePxO9O95bzOiMrEG8yhHKerGXf9/SdXoKb8PbFP58VvGbEXA9f00T02w
ClkctjPGwl3s6YBOGQ5nayTiEUvmQoiWZdUbXVUwwqO0XqwrWKIateiPLij9od8k
lNspJJ4yqmmQlcXTSsYtXS5oBDMQ7Rh9nleZ9l3ZK714clz+KtKcK7kehhA8ugR5
hsQ0VIdrCVhWGfM5hvjtyMgJh3tjv6u+r5+q/FYruMEZLFKDD5Fxb0NX6+uJqksN
+BlLS+q94xxqAK1IUWB87hqnSfZcGR/N5mpRQCzYC2WN78PxN4jfxyj1FSMOGK7z
UDvzb4x6lj5zeTBGLwY68GBgXww0k8wkzqACzSMShkdNtpzmRSlVIjdyfjMO04PZ
/bNp0ZL5v/qm76Zl5v59i8BAGG7ZV7zhsZHgbD0O/OAmUkDga4eDQmRsgfElF0cJ
M+hN4EuaYYXVx7aNUO99p/xOHiJ0Wb87nDuTzttN4PqUVv+L/v1jdIU3edYtpIYe
LkPYNWieX6qAP6ILLzZBgtaJg8pTKhDnC2756xaMpYjmSDG7Uboz5ULUP/9WLvbv
SP/l5z7Vlgu+ewM/P3P68xbyH+Wnk52viDSoJdm4sy+pQ6ofoPdWioPXr+1tO7Fo
TKv6uZZbNTpb2AYuga5XD9/eM3zBMNzCy3J7Sfs8Key7KQSJNp+/6Gc/qfm910Du
M/TigzGOn66EJZRMjFuuSVd3JW0h5RIAmh4Z60cI/3HgxPg/fWzq81Z8Chr5efQb
doSKaSVuendgFbsuRlO+lYQFPirLBXleaOzzP+tOp7FSdKKxAj7szG8wpr09as+/
c3IZ3SDIbOjdGNdkPCk1oVv+QzYLsZ4d6meBlsR27QQjp9YObLCv+8L8GjnqFStZ
1SjXfi7+dr1Nq+Y5PGe4B2PhY1KHJmaP5rqoGiHZUoZYsUpc234QJFi7aUFrnR+W
JtLkbmpqd6xGUNntaFCu3lDKht9792kJnQHcys/PbOuDSi07JWRZkSX2k59YHN4c
f4PBmdgDRPzXJFTgVED6E3hAGmFaNA3+Y7oVXshkf+ksJKcONr163ZV5vB4TeFyl
+7f4hvWXDLTSpXMsc5pYA/PhQXtu8zdZskkT1QRzIezrn+q+64Vg2hR25ODM7ak+
XOKLZTGiePXzJp/ekuIlhVl02GRfUBtXG7pN4atzCo2RB3AQggoO1Nr1HiHXv3sW
E9XoKdNi+OiIV91KqmliAilRn4sNelKDTtzyL/beBy5LN3at8VkNtFj84QIbv3pE
cF0X1Byoho1W1JiEJDK9YyKcPsNEPLHb47sToSI5kX380wgDYPtbrwcZIt8AJYHG
cBIeJiNVphlsUR6f+KHMyC0IRNnerhpgIjYClC7W10t66bAfNYVn1I178tnIfouM
TaIUPiK3+qFuy9zyalHbE3Bkup9jTRptNbyp5DmhTaHxHnrh18JKP7rGldjXFQWZ
sViEX46cfEClLP696Cc+cj7Q0XgcCuEYPCvH5l9jGkDebI0srNvyYLX4wu7rXjhT
OFU6S9QGFwDo1x3VtmhWMTZ5Fa43TBJj1bCfJG1qEVbCV36D7BSEVSdc066UUN5s
zOmIEbjvgyDPYqCGGuSKLNyZ/e5zSYkyMFc836vnvDG6WciOGmPFF776ESBBfQ3e
EmF8pA0b9UX6D7opgU2L3Cua3R3qlYmMsqCcS7YIFWdX8PkdOWepRz2UOxDUljis
ybdMH8v9UUKbI7yStvDrAxz20gnIvrYvvyIrl/nW5ZEngML+nFt/0NJyk29ZPlZ1
RooWuWrwtx1rlDIk+DxEvWjTD1xp3Rg0pW/obvl+muVDN6+ppsbkTHG/uSrXgund
XAaEgHAXO4WD4Gbg/lELzPjxRtdQQwDN8SflIMajPoMg5tKw+qKhwN0D+AFXODiy
oEU0Zg+aN31Qo2TRTBvEaVLlTo0IjnsciDGZkRNI334vb54IWI+Kh5XDLaRRWVqI
qPkIsMT8ANqX9yG5Pq5tp5Xo3D/QfeHRDSw7A96PtdGnmD1XmojCLxqUj2jND1qu
v+Kh+3C/UmZcmAKBqNKEYRGlyA4OWjBhxMkz90mhpkvU6vYEwR0XwbazuuBFBZeo
Tr5dBmvfN2hFy0PVE/RuR+wF7sLtJO7wGlJYOXMnntNQ8t3MsZhVF6c3Pm2DwIIk
U5CJqEhXEgSPQFWtzzrNiabdhhcgaBxcVYfjch50HJx/Hq7AmfZ2W37GU6ErJRjg
BiTFbudAXEcrTN+tFUMrByo3fZdW55mjPyGbpbXXix1uWU85c5xTT9xiqCRZUcfn
QsdO/waCyLFo9xp4Iy5Y9VHKDDyabJgIhzZyPudVFp1ajta6gXU5JgA0R9DujGdE
/5jssZ5wpFSi/pZGP5aPl5l5vxFrY8va6BioAS/KCjy11reEQotZlWsbCdPgrMzt
VgNy4E4HPzhJostOKTVZns7G6TAllGBto2px8ZmFqlgpZSdKe+x75vj9NlQnGOBZ
TPPBlOyjE6z2zFpC/PKENzzDUtA0RfKt7ogVZ9rHaeEYP5YiNaNZBSp+02VSaOrm
Xzu4V0KhPu7ufCZbXWStaMjBtAl4Mr4CyqUhHPIqYRh+FTgauY+feY5pcTySk2A7
VZ8onE9rmscCttYhSRlr8XkCFJRes5i/dPD/lFI4e9Ttc9P3qqchRoI8ngSFNKFC
ZoYuvtkKEadmBomWIonFpVqk1bq6qIScRZAis78ddhh0TomDBoHQKUOXvlCP9rgo
tWFirnVVUMxPO39ZsBBf96tM0sYVJ70H/GTkAeVfxMcyKLJjNopynfH1l9Un89VB
MddqkBrqMvS76LQS9TQwJwQ+q0WE2xyZ57GCF9p6uhL2yIpar7f1dR+47A+39hq1
jExfBeh8V164zMy6N8ROev+2bRO3lKS2+ULiHluPtPg0f1O+VkuYdMqAewlWDyVo
/1DlL93tofRSB/1fY6V5SScmU5fM6fImiUl9n3ISzOf2HdsjrAcTmOHWvRpAIx9a
iWRorrTazFVuiiGaCQHdRSvCW5d+TLE2q+rf6EElKKVPwyolHU1FTW238eLYx+0P
wn6FZvWY2ys+OXWhTVbAvdjmwjOfEIfebvfjZkLTF8l63xhZnfzZioQOEDlzvHwY
L8xtehQBbgpR8LQZfTVwIFXxK2+PMxeXwsdR5+tvvEcB2x5pasD2AM/KOswDL92a
QdX3+L4WaBCPn+oG580naNzhzg0zZyandzP52hNJ8mdaUn+bmZmNLWhn4sl868lP
xFA1zMRvNMGOhgKuyLUKsbfGoKJrZm5ng3fOTN6GKmjQ4YM/pWJCz6s6NEAJWvB5
N0xR/ZpL1CnmeAQD7OwglqIYuq+T3DYtrw+kVlLO/frDjgb1VwPu19lEkMODHVzK
Jueb57ACQ1JcFjQqU0HJFEQjxOU4oqfWygfZnDbo4Ss4vgKVsQYQwVKeMT9URe7P
xZADq/rgDA7crO75F0XYipSIgh7MjhqT2oCujjGto+hFbV5bcJWvLgxxXeKRQ5JW
+g3G5rEN4qSLr9E9cbvcpeXERFxZ8QeXoZrd+pKBRbEaJqBl+HORu6xcAH6Z4Sgq
AHB4plg/oqFRLvqL66r+UNx6wCp5Qa80ujNK1ZQEDLRvyX98pVX2jOGRbEAj6oHB
8/r0DwRtOu++ibcaYJA6Wevo7CcDqAY/qvhMPbhfTpDUb7SxkApYhCIKWKVJphv6
8ZyWPEBBNSIui2pwAAY8HDBZ/9NMOaRhM2vbp2kVg/R/DRg+oxITWkOAPu2DVQcx
GoQ3JqgJEw35E8WcI1GvAKMgl7gHIEJf91uNFi1T9hbhaqmOkSRswbwiJCcCq33g
tO6gvOmygmvdyPudJIY+WcYijTyf3BL5NyMVbLK7lvgij17iZt6aHnb2WBZE8ud0
gFemg/49VOzm/xOrd7S9SGT9xgxUGVrN8cUEWsUcicsgiCrb+nA8GBUyZgaO5u+l
Gm/cybPlAx4ZHFm6ACKEw8tp6IVUMwdsmktVqe1l+v7gHsODD/NDELZCyfIShzPh
AknjwzSMp4wriScm1xtB7v9dkQLODnPItNc8iY1MVggualC/4j+Cc2M84qI8MWXM
KFiPvZujXCyFfBrDLtIfkgWYN/EhUVGUJj68pF6F4kDtCy3NuuCYz3D2Ts6BzC/Y
EODc9IE3RkoZP1W3WG+F2zy3s+HtXMg+RVc9d7B5dFsmgJhPR3/P1PMSV+Z0IWfv
ppQQfclzF9EC76/FC4ydFg0Ezk3iJt3imf8fJHlUte3EB6qKYGMH82wRtMb6XQEA
/c4uplZwPrln3noe9i/4YqN/GtIrfOg1kWQCAUt3P+21zzW+Q/axITI8ycNQMoEW
NQpy9lR+2RsGSTodij35RkU272AAhGyu5TlILldp0J0+iWJvDpg4m/NNq557c0TL
unNJxyHxQm08wxOgYYHajeJEr1xlXXzQIfu6MfULdEgwLbjQpq543/+0F/Z5RFqX
jidv2QvjoXOZLvN4DMP1uKpYoPT70+nI8C5vNB+X/kLwPVYvPqLgbGzUjRSbjaJ6
BqadNj9NVWvlyQcz/R1oquqTEjqM0W1bdm0HyRQ/fFHbWlZjJi5Ec+9TTBw+6tw0
nHrbOJPbpvtXEcIw6I4KFPpQPFVbP0Q6TB3S6v7YSY0YHSiCrVxCiv6CAGV3xDDj
ryTtTgSb+lTx2nCg4ANt4X52YCVlTPrV98+Sd6Fo6QIZHrUROsJShaabGvHoRi7c
JUGCDUF2f+pfLP20QieYbrf/r45oN0BaPQ/fut2W5zVtwrCGfD0KwdtXY00N3liF
GVhZNoUszL9Bdl6ukOxe4g6/sA9HOQ73nW4IH3P9FIxRH6wVkG3AtZO7Gg1L1Prj
5Qe+zLvp5l/H2sC+6spdhq35lM6MkQDzrObgzVmjqEGcvBcUE4qW3UO54uhip2cO
vMamEw+h+MLnWX2MLClL1aLhe47L8VHKrkQKP0kGSs67r5q9vBXB8ynPxuy463q8
vMfYteYF4zjrcFxAHeoYFrQxKMpG2t88o8s9BTOhNL33e9Ew4KGaRhZXreGC3phd
fRUterP/dSKd62AcqrWgclgi3SWGrQjotVS7mK0aW1NtXDkXQlhP/kvHfJSbhTSN
e03zY1T9AvD9kYcGf7aGfC6KVbg1doQLeiVtqhwPvxBIrCRIrxnNC4mkj4NAdd3e
zILG7rUaLGKbP/oIX44g/dYQu4NHDq2e8/oQn89IoLaKeHOGuN6JPlKybjxEHOvD
YFkNAU5ZE9t8iYizi2MOM7XsXpp/C8Tn+nZWp0XOkwHxsZflpRPIE6I0i/tzXY8w
PgCy2YFh9jgpZQunQ9qy6vWVkjEUMbrO3ME8STPVPjIA8uXMNY/43l5nsNMfl1Zr
7g/+QA8gkOY5GcRpYoFVbnnsxIQ1OLobAhp7GM2NNoHi2wURMzlcIiDta8UgttS/
qTlK9n0BScwYO4E5fpIHI25UCUQrkVBOTNbtl/Dy9p0c5+KLd2Wgkfy9i8GwG3Uo
sAzloZi6IDagigZEItvZlnJA2aBGfIg6bg4KjeS6ItFFX2NJnTN6WOk4rlOnJtQf
yBcSXicbDmDXlakaFt4zOZT9NwDuAKTnuCD3r3Qek2QnFOVFN43wNym33EQZj74I
MalqzIn32jMkdmW8QjAeO6KdPcN/h+by5vAThEh3X9PUJ9GLiSHA6QzMBjPqLW7Y
QANS7ltfFpJVVe3dzH5CvlE5/X+ExtAEAgUOlPs69mpXHJHBIda47Llylp1wADwW
pfDIXoIidumCJsv1mbvB3ulVzikCIDU+vw+ltZ/MIvOHHeWVhvWQ/y4lq8sBpbKP
qSzGqtH3r2zIn+BDxBFdes/V4Xb4Z+jB/YemFSPubkroH/vjJh+etDR2pnrUpeHk
W+EqSRbBnrpscwU2aNDM3HbleYTde084vh2kvZvjCgnmFXKZMTwMTv0uwMlkpb1b
MSlH++2c7nST+kMTca3AffkOo0v44UMhN/zXA/mtTbgjZtZGXnUUY8p0xLi7WPCm
ncldl/CkYLC9Fe4sM4zgeKniD/YA07tF9BlTRYpHcYJ9ZA7MK3Dc+p1NOEAavelX
wsmzpq+2oxU0FWFKzdqQjImK9lXlII7yekXB4ZoqKuj7u+8/zm6PSBJAncEj38IM
hCKTu2lFTrQ6dM7zdvyDys2xj1wJ9Sl9pploruDB2Lll7fgjSOCGLApk8+ZvzfzJ
DDjhcYrBEt1Ms33bwgwe/bZ2jPQjAXrCA+AJ4jE28piCvj9b7VA4uX+cf5FRTwEc
QCyuKY2DJFMu0/2qk8rHbdp2nkmxEjfwY60tPw3LNyWsfLdHzJgz5XGzKEU36qG3
ilcC0i7M8RA3FGgx5eBrjnaLXwFYRHOVgIZDKVAzX/85X6utsJ5XgYwfNuz9w0jE
Kn1XR5tGoKKiMRFH1s+w2COSUuWnpQfG/5Lp33BZbjUPDHi3FOG7ftmE+eeF7njF
5uwB+HJ5neCJmkgI1RlPTOHutWMMEmlbNPBj6+uDVZ6fkFVukNbDe9iCgQMTibD2
kqNrp9NgZFSI2cN34pm83RpwspW99nmCUBEE5sCXn+1/XUBQRazuselARsTCQCQN
y5ObqsmoQJpLReBh6muCiIP/XFUitKQ+KpUMQeuO3OzEIHb08aNwobbFDinfpwBR
mKoMOqpG1Tj1lt9y/3R3sSER9NInukB+Xbdzh6km8xu5fDVb7hYbINgsWUamLG9A
V1ThEoiH9vmy2jqbeCQ18gmJA7zdpg+w3qg+HlBVEwzy+ObmPH0F1HAvKbdNA37f
Au7amQCk368YCY149yaMqMo0tqb0lr7adT+EYK2k60o8KLn89P/p8tk8bETScBnz
Gs8OamfTqNZHI3k++cK4b78VqYFmltzTSlcGsHomW3SG0q4wBORle657jPlryyEI
w8TYB4N3dyHDU35tWiwvk7/PQiwvduRvpTGhoNFSg+eyH+6DPt8doOytL2bF+34f
y4s7pQaWlgM4cERFmR6dZLCPmEBVe/D2jbSP4Yn1v9ttLYDTruk9sPKpbMMNtpRX
0MdcFKg898r8m1BwkZykN2hrdvnEtTUzrcRl5+Qh/MB6hXNsulX0UNaaGr1G5THz
7oYLLkz1fcvHJhZ1qeIaumiedxSQqHT7VQ8DH3nbKaz0NZd58ity//M1/MBfEjDM
nYvR22inXQM7lrWeqaQn7P50mkT6OFJ+bRu3vsurpv9M8ui8ppbptzAdh/T8uOD1
5rHb5bbhiHEfur0uR+wnzNAMhrNOJHqz31xp+ldeevcsVa+H0Xgg5QCMXFIoNIpy
DFGyexUUV026lO2Yusm+9pW3E7iplc3NQtU4efbQcUeRFmE2ukSXuTRaGYUEq6Al
qEAB1cdNbf2sBb9Glzyyt5huNW2STT7fahs1Zl3w3zjonymN2EalzXVc3uTH9WBL
B0ga8Oi37NSUWK8vbeXZKp9U5hg8EJfgoO3pCk47MAi/krhaMI9L7nTA4E/tbP9x
biLM+/PEyLPYjv2l8xFzoEY8QheX5fApKis5Ss/iAtYBpkKihRkrUKsnyXbYzszM
Fs+88NUz6HVCjVJSxqjO0eXiZbXVh2CKI3jHbIYTsgbP8eWJcN7CgEkUoxfw326J
LZIK6Koens+cowiZCYEaITEpz7UFCehUqIRt7DWvm3XhamA6miFUXgh9YaMuPqos
8fXUdv7T2cDVeUtu5l8exvIz5gwYdqS90OdEDo64rrD+xM8QYW0fC5S3ZeGmZyQ3
LSBfuFgw9wM8Jkt1rkM6lgng+6EK/J5AwGa0hEwtHfwHmTfY1hq+MpAKq7N5Q5Vu
Tf58nU+DbQ0Qi7j5uAA0u010QeTllxMgHd0XiBkMIwXJczFNnkmDWr7dmaQnfSWq
zjKnOTHULNqfH6LV2+iFr1zbEv9Xz0R5Tk5pj2WTfhhMuQFnbDlCDRODv6Yk+VkZ
o2zPa6PHQCb5l4OGK9Lhp/FYd7lVRQwLh2hhNeAbjNxjglHm/ArSg9wFLLw7FR9k
pJMe2MdbxbnnCxUSLGtxGfHFXXIoihsw3gN5UlZqPOod9wfkSBngMlz0hLkuKknU
dmlLLTRJCywluRkDOzC+8FmXwHMj660fmH/85gzfIYSxZWPXV/I2NJ+FRR7XJOXA
Irn9LtHIkvOueCmHgfUvPuQwBbqKYIaKvhJ41DmPlDsX6ni0mLP2qPx24tfzIDKM
b2adLEjRH+qiw/c78ZVaN51FoSz6fNWQ4tfbrcWteLlFNGKJ060bJit6zcBgEP4X
i5Fdbm/13pWByvZd4+i8U6zqZ73Df/ysApgCerb//zqeozIk+9CjdnUwlbsDDZYM
8Af1zrgTVFhzqN7/4mTrBQr/bMb2jp5g9EErmijvoQkn7NhikYc7Q6ok7C7AjQOk
ZxmBp5IoZSJrwMC1Px7rWudY9MQjh0xJwoCmTgb6vxjLuuqxZyKWUtQWL8spccC1
/2muAgkjAclU3Xw+ay9uZkciicgNm28CJkId7u1WCLW+wpI+2hfCNfsQmX9YPdXz
yuP6gt5zMSI20yKO0mFRt+z0XCydT01VSqdHejOXN4VhpGJrazCj0Xq0tkTQ+6HO
ERF33XM/qnmDapGS+N7Ga9qtrfGBy+ZEkyfgoKx2j7K1Oj62LBHx98l/3HqVxokw
024vj8s3eVGF0SzzOXqzeaF4OqkXUCPwJxQ0+EMDWjDcW4YxG05GO15J0m4mL/Vf
sHaHZa5VZkH8DFiKKJd1Uq7HvJSXk5bQv7uPqj8yYH4qFP6xc4VCwuM7/SOBgHUV
3MJSXAXcZMbhsPFHKK08lhp/HepJ1oFX7Jjg0LCyVoonfDJUmf562gpay9QOPk8r
I4IzQIt90/L8KGsh+558csWeXgL5U0P1wvpZRnyYrjaXDHZmin0E/Wz0u6aypcvi
ZDyef1bdh/fYytoU3T0ljncJPjtYx8JuA+VeMa0xHU29HN5x/vYQqgLcw9nqtelw
qXHWqWq6zI26qDFZ4JKoqJ8ohSFkJ1WJ9SLE65HOf98m0c9p1WT2NmonSgYC2RIz
4as5abTUTwgewyXfZbM/EuTwf4audbHb55O+wPPazGZ5M0qML2pB/+08aVrmO+b4
w25GP0n4EqDt30ogL1j901yZ1j6zz/TmpHhK46fYKlooadHfALJMUeujwDXYGVeV
Gisw1glpTy2Qb7f23Fr8QezZ/wxcEAQ13MF06ccg7a7gfMvRtpIjjkG+Sl6NEYvy
M7NFoupn577G3j+fSWbK8xtpXIpEUUDRGaG+mlQDEPtOzo5JayJOOJz4TGwphHc7
SGCy1eJtLNfLy94i/9NF7xdjJ7Iojirn7ZEFIVTVpY+3c2yFXhZGQFSoUs2jFjUv
MdUSYPA/w5k9tysPQJpzHK6SBHx+JfXaJXhXV7qiwgvNaNUhGp0pP8vO7woR2zrU
ho2BjHvdk5WqpEHVLs9WxzWF+D4tMpvMv+ezughT/hoa7WXnCF9ypycOONnV8V4s
ecgDKS1VPVtt4UBGWpPjybJnUiphqnEjcpS15pzK1PgNCAmBRZMHnNLjLN5GsxlO
BH1vkCKzo1dpXuMyT+LHZlSqZdVS3XdlpdSP0ji4VtX1lZGNJV7FS/zZOWvo3zod
NFWYxPUE847mLGYi7pG/0Je9+xIXWr4ziuEkXW1IXI9BZWNVL9svka/xSA3CBmvf
yR5AoYtHtxpZjmaYqy9HJLk8oEFqR9nSf4ZGXBz3lrIH0jnKluO4FpBqIVcrqNRX
cy8yNXrpsJp/SX5R17IKPaP1PA/OA/srx7T6ekWJKXUTYV+j8csA0eM310UhsLwg
zpI0hxiqrf+PAvbkyYXxoxalUBXFQ2aJ30Mih9uXqWwSE6itXM4CkJmqhpg9V5eF
4+BtM1jGH3bUmrlYBxEewjWY1IKc8QfC4XoIabDZNAMVzJ8xp/3okTbR7/AgNS3P
g00v2Eh7OuvBhjgNflyBRJI7rB2WOoLhbVEd8bOTQPnSJCJnSa5BQcbA/zLmflhM
LQuKYyQHjFSPxeqVPhzYKO13UFGKXlHzj5PisD6YKNWQqBm0MFYMooGoguU0jgu7
LC4KklNJPI2c/VZnEq3Y9K51V/J43w3p44iskCGd5nzsIuKNxoMdb21cphNzi3Pn
g27wJNQIjFI4usvBcPXSHMk4DBRSUS9L5y11CjuxN0s4GzcqtA/sxUEU4grlzYXO
oXW+WV0ImKCk8eG+nePWxyZmHX+E6beQzW0KJ6TspWXcWmlu35P3xqNCcvEA1j8I
mKj6xiz8uGuwqOivIBvR7a4Vw8TUB6S3J0uYOF5RNPDpYarW101HPUT9eRLBXbsp
x6SXXnbNKvBr+IvsadPgr3BIwAEEN7plL1MKR2AQtWk8AFIeoXxg6JIcJFnqRmBC
J7WdHBWfhhADpN1p4QLLguBwTrhflfw5ZpZrgaYLcCIQ1NRtB1r4zSHHvvW71zEF
iLZf4zf+Be0CUzbX+Uq+tfhseFfd0cSTyVHoWJNKz7R+TI/qeLKua6CdPcqkhrry
pbMywr+I0kiMh5PMCnIBO3Ut7OqLX10ClaMF4yTiYgBk70pWcQ+l8Yl8H7lInGA8
TQemfHNSIxSJOxbPvfF4F+sVh0HIBQcmlDueO2XOdJizuL2dhLeVGyBE0G1AQSXp
2Wdt663ZpmNNpKgynw7UREHVazs0ySeFTlg4IY/nhTbrenwQ6nAMxgycmwguGPiP
j5qSy5tEFkpa8lag9BPEgERFGs5LCORDgKlFgk0uL2i4xSMcaaVjtzboLJDZCh7K
4WzzlVPKUsyiORp+gCAmPp6dToZJkfpSP6HLyIRM/LYPHTeKu0T/02vLGaS+Cjei
kZ45Zkvkt1k/th59fUqRve5sBo24NeKyW+FGSZR07asqHEvPHV8KNYWIB4UPp/ds
GbG8J4KUDkl9upmo8dVusD29NR4V80sWHt/4c91fMNPO9huemtnA3vBE2kQhLsJX
HKA+jBcEexb0RdQBZBU3FZQFAz6Y3lFHBNZovPrIsDv7xu/n+QIV+AReEERxrmd+
eTHtf/kFmXMiYwfJKCFdKBxwtcopZEe67NfsOpaZzL3JTenYccDNNqbiZgF1umDr
Vf/Rt1Fze+VtTAdUTS5GUJL048FvOFrZEPFqHYgOfSu7YnyWbxK7YywJEUVPrwgT
fgIBSIcIYJeFsWlHyv6Trv1tJgPFuqtcQVsKMUfRzvUXyU9eawiHFeCbyi4fwYVY
fYmzPhtjIFDO6fP2kDGXcyUt3Kf7hi07aQejXzM1pOxBzoekfCpqOrcR7PJU4DFI
bbYP7gZPwTcu88YTJ8AOeVWoCuoXB+vvxFkqE94+WQxpgSTiYyyV1E7NatKTTSAV
/81gykC2PX80Ox/PM+mbK8DCfV62FHz1z+ohi523GLSRO+ZZy7WwYxL6dRbVOTfl
iJPduxGTwG7uo/LWpDG7L/0duacsbp07q8HfQHtFjdCdlWJfXHedO38QQrd9g3jL
mhJMvwjtP2S/c3ZOyopJDuLtb92qEryMJI6zoGzWZqyjoT56le+6Aqp6rNn7Wa1G
7X1JmbYiKDmvylo5+ej28I3/J5qeL7Zu161Qais6zXutRWfTm95fOkp7nDIjwXe2
P3QnNZ4kQhrPOUIDtW1maHnKxuHmgw+Au/eAeo3onMUcO8DO3Kvtkaszvb9LxV05
MO5DcH3iz/kpfmLOkApEK9K64mOhDOh5XDt4AEkrU8IY9WfEyJ5lQvoDH6KAsxPM
wxXZ8Jglr0twRAx25ubvcQANk9ewwy2TMj77FatZdkEUEfS3swSOBCo5ob/gXGF1
WzsEsQlaSa5z8Fkc1xSoGar4/XWerKqvsXZQ/OU1zLhpHv+Bgrgg72+TThCpjN4d
C79zxTOzIgC8mep/X9mKm/GStl1wrVy77aogGsm8WIZ6fEDGwSZvkz09KDYLC5Gs
tD1iOi/7ZEcm4q5qmLRn+dkWgp6+HTdOCeVA2vpRo8TrIX7zl5p6mekz2wN19TCq
FDF+l4uvo5mG3hMY/s0R4bL7F+Rsw+KZkLYvptBLI+OgbDVnQfqPN7DF2MhVY0Ui
YPUhhdoaFIu02b++QGsjv5AbAQo+Dyjaq2toEIygDdD9Gtjl8c0oAyIC25bADD8A
mYXKmfIYkiXf2irevSEcgeyt7OQ/aEEEdpXZEGaQ2lEa7FOVvSalwIdgPPyhqV7a
wGIMO1QoHluC1HJ3AOcCoMD1vGq4xEQUPMm4UpFR55mIhB7oRn2ASbVnHbRx9uLg
V55jWTDxMq0jbglc1pS7eoyPzEUHqXUNl62p0Ofda7bWQ41B/jqCdSatuooE/pJh
3YDieKwPUyhH6skocfPd1gwBOTjm2eJ0KXFJtpkLzgo1IejUuIj0ZZovAF2ItJ+5
ERCYERPrAL+bZUZqcUx0GnoPef9C+V07OBjD3WagFTRvnn+63fFrNQD4GUdUNEBz
o9Foi6ARYMly+uUvd66FAXID1yEJFTHcvNfTJ5ISBhB0ZmHEBkXu97Rkb3OWemgR
3iRr1tCLm0Qdu2oSaGjxyjYdIhQbGztoGjc0iY9IbhQV8QWnJRNBGAR8qlQkOaZc
a6KAgJdXF+dDnlTlDIy2vAU5VNnx+qxVGibBIu0nFn5yupU8wXRyFCeBRC69PXKk
xQOXTYTa1bKN3CySLiBokisGe55Vs08nL5Wg/HpVtrILPA/leN0muK/uvgyiV2v5
yveMrXRoMVW6qwa9CNbbLFnVFS3SoQ47sD2O4hUTMzRtjOeb8HQuvZi4A0AmLd9u
IOeOIleoqoEFAgZy0JYcHAjzfCG9e9b3nOIRwAHr2wBYS2DPC5oYAm44gyPZL6T0
lNlIbVVDO/248OYgu8sqvkjsrZHtpj/1hx1fD7gakSaamiKyrME7tmdHHtA+BD+d
guhksTEm1Y7tTJVj8PscwKiDkCPfYDWX/sjJQozsCajC6j0xYbs3rJa9rFWAmUmy
FsWiY0EMFRAk47qFrDpF3cnyiHwDvkbSxdJNspz8vYSWQsl7JzUx2/5VqSdubhnM
B4PY/Xf3iCcPybU82r1xDkH6YnX8colKNfRNhYJJ4JpbldfqZQIRTktpiTbNRq/1
Ls2M2EraHKtgWIL1ENS6DZFpAwQgy5HBP8ZCGgYD1LV70gt2w3zgxxawlu8IUTuL
Y907AOEwTFHMlrNAekW2FIYc+gqSHQWvBOOE/Vh1fqEzCpdjbP7ka3COD3JZkpbG
XqnKmOLAUIUzhy7gzGTuqvQsUldcqxe/3RcvGONY6ndFnxOiOVAshfv4yIe4qo4+
J9g43gYS0LHkjaW52BLbCFTImgNQz9BZc0ZovEeB1vd1iU41SwPaoKRrpE3WMlkr
47KFYDNfvKx7P48d7UId/DFmLOoentgrQFp/XtG669IAyReZA5jLS8vdJAQCX+gl
fCYalY5sgE5IQCZSIQX7ULMzYZi7stkZz3dLPoDxwv1u80C2YhfgOkxnx9Yc1oig
Yp4ub5OVTw6mWadISX9lJnqTfX1YkFGfwJ4F4RlVM5CDJy2xq0PKjl2Oa22UP8+b
/Gh/oHGDN55JufLA+kokHrNett4EvYesVkNZAVc/s55QJW85RrMy/sEdZWwR/9L5
J3yK7lnx81j+EVN8P++O1TIjmoyz0pgzOua1SJK3SKx1xm56wm5NxMlQzJ6B11+X
/CeBgiU6bxnumjRljYqnVww8DXd8eaYxNSYjiSH8j/1QBoC7WDakzIDgzkblsc5F
PuHIjeaRd3zDE6kEB13KGLQquM4r0vVeh4LwrFW6fiMm64KJnCstdLYgG5HZ7UKx
GbmGLCuggOGUztPKvVgHXhuryPHjiB0F0uw52f2y+uWJTnT4ET5aHv6pwcEEwsOs
uMRxDE06FbDQSe70S7Tk3X7m1CuzYsMXhLjW/u2+B5PaFVCGq7wPeGYxyzrTISPw
TuOFQlIxYDLL/hcm5ZDSZjg6xPRaAo5rvf8n6Eghf0UUZnLPrp+GpneMJBojV71I
eSStOTk03IVTwo1fEtui+W+u8XVnuUXfzbwIiS2FLkG35XlyOavAQzGsqXOsxICy
wi5OZCQgcQO8HmX6m6I7hals43CM2LZsT/qP5gebaChxuJRMVzZ6hY4HNp8pfe+B
RvGBtGiKKX28LsmjIlydUFhADwKDWwk/eax89jjBH+XPHCxSmTUHlZlhxK+HijwN
EWS45GwNhAKxB1a4y5vKM43aC1M/c5ANagrPr8VZTWsCqeXQfPbP9Ly8ejsBuLmK
xlq8RSoohs96rgfxH+R2ygvg4UGJMpZMpF99sZY77wHJrM+wOHo0CVF52fC92lWA
0OKYgOW+1iqgTckekI54jYfnrhZAwY3kiCbrvkXSsag7Z1/HsZvKr4X0UrINg98i
9/zqxJkn1HATE7TizpypnBv+92gMybaIaCqS+unKhaGlVu+KKrTxmlt5zzZuWQLc
QZTm0xqRC0+JYsO6A5/6Fj9Egtyyn2CLBJlDY46gq84FwgwfLUlzjT6/NDZay/FG
BxRISj/9HGyNjxCEgF6F5dMxAJnNxR+1GQ0FtGuc7ZYtU9q3s/KoZMTgx3XIJgnc
kRtZb9JRiEA4YVsIB+RA3ztHe3wgck/Bok47fepmMmu5kY+RLvBFah4iZLLtzEt8
bd9XbSZvJ0rNKHnpri/ci9a42EXim3t7SXgfvcbptv6i3ogbaRltMFVXhhtcYH6R
FeOB3lDSrDqZA+jGj1lXhxzr0XBahOIyO/Q5S7yhtbDgzil9KpxkiIn/5wBuk1Oe
/RoX2xlavZXRa0g9MWKXiwU/74z0UcYd2xdLbmiRFEHs2sNkv6R32SbASRp7iBTg
b2gV5ShYvDHcKUAoEen3UUJBzen1MNtFjKx+Hy8tqKDUnhuOjsc6hRkPIAyfSg8H
7vYl7Sriirt7gnqHP1f19JhysiQQ0aVYsvxkoLIhmNdXGUzQRix++jeDSfeBJTk8
jhOJI7Gndu6sRoUy+sPAhQWeyU7cDn4p2QX95mEwHnzK1oSoC+tU/B/tXJhETbei
eO0PLE/tF6RQuTUI8dkXDB8WpJUwn3/LNLauLRw2IzNDfUEXrB2v9kXfXurj7RCR
tdG/aL5a/8r2HmkirgFQgebhe9Vra+Nwtr0sT1usj/i0UbQM3HWLHVUddDqhzaEy
RnWOdtCsLkkRUjps02/GYWqCgJ6yfbvmPQXWQ0MuUK8rDGMH8VjYYU71wTaB9EIE
qRYoo2J9Fd0lqj4CuRcJ7PgakdcAUiBH1XVllQffuHRYQe9xao67OIo5/6DuR5mI
+OQCFDWrITOqB46Dm8+MZUNiCJ503ZafrSlSDPhluN7znkJBoF5b9rdf1le/zZEp
9V0OOrc+wdKx7xbpyVN+3aTJVQzKcpQ4ULV40GhH/6iINlYtShWRMqc3wNQzNW/6
LxzSAMqDxVkPs+cCTsxwvDbMrL5ixiCCukKZs6oDiHg8lMcYB2gqgFY5bIcu/AyC
F+A8gwceGTRiOeTdPwca1axDdoDK/wPzd0OudCU33Ovp2f2hI+Ny3jrvpwSsmnaf
+Y+a2mIT11dXFoh3vTVVrLqirSl1DvuVN0exqJlSm6NUSLscZZqsRYFllL7qHt9i
fGXljYMHEDOj6P/Y2kxprcii4OalsmfEnZAdyBl8gLfLLIE3RCrlLHQYgh1Qp3sh
K72zQk4utw67eNhbWertxFDVqzCXFv1NpXfIapzIrPmkfupjBd9+Pe/o4xk9Xqvx
7mMDYcMs9zDvh9R6YauLkb7FiUW+PGQx/mYM/JcUczU2DPOaWnJfQWaanuhzl7Rb
A6U2Y3bUW4lnp45V3SZr40hMKU+4l7ZHqw9M3sW4p+S25Mmyy4kf7LDaO/r1N7Vx
ezxkp84d+E07N5bTkw0vJ6pEamczE7aOMWJJ0xxU0Pj1Uu74FFQZGE/AOBoEirAc
/X7ZWs2IKfxKD/7qPDrJV/bMz/eQEaUVyKen3LZK0FBcO49pK6IeGJhDnvORugoC
HJNFNLvUCyb4miBpjdcm7nliCMxbvh8nDlw7sSMyivgWlzD9WQupnDqamMfYqGB4
LSg23wzsF7AobvTWI+2+5QrLav/UxwOp0JGEmOuUDGvomicfGpPtN1V/31MgeDvV
WupzwYT0uCIOArcDgbFualpgte6UThGfz/HPRTn6QgAF5IH4l1Jq5R79Brl+hoh7
MPpKN1IzhTrLCjGKfapgubb43494TiQ4oLknF9GI+5pAu5ARMP1fP3CYcf174htp
iy+nAb41Ws1ow1EAodZasZYykRZ7aUia4NBa4V0P5z+DsHHS119lZLhZBkx100Ff
2h/JhBdZhai7iZuWG+TuGfpFvWSP7VBV0YWfQ82XRhn7AFdUR49GWqjwkAzU9TPI
o7nFecQUcvTlhN6Ctk0Z8GdHbe6uZNAJALpGLPoMlxvLrpQOxw8MySl2aUHSUxPg
kSvCzB1M02jwXwHD+kG4Cubo9SwmwOj0sW5cAnzU0hK/vAi9iu0ku7RCFptGnlCA
0VJUfv2SBQl9Peb9TUc8NWd0WCN7+AtdWYidepBxhq+ZaSjtWUHmi3VhnzBGjCy/
iaNmP3EhnSm5tbSZ4z+o60ZKVoV2LxViSjtF5FsiUJJIO6KogepPSFPaZdOnN5YN
5moyk1Ph84sNMabDmf+H/SQ2XkzmJXBRdaiBNQQ1VvvtySKJ5uD7Hj4eIyIrUFbm
IzVrGI6MNo64E28e8sV1vPNt0Dg0P2TCBsnL4qaYajURRwOADWoRXFjiYGD+HNkh
aLVxCo23t6+02eDig9fIWGe1/Wxe0/OLx+Rsjcj3zKSv+jG1o5qpJ9gAtpKWqnXp
CjoajhTnPTJadPfgEXXzu2u/2gDPFLXdn/YN5Gs2v/fufjy5RIwd2b8AvjVo2lMa
QhHZiILibSqeGl9zc3rf5iYUQFXV/83biPIPdrdwzWVALNyGbd/jnavd61BLKh0E
r7NcmNG+1XUI8RdvWJ/0qLJezoBMVp0H1nfimNLVWEmUOeY0oHg+y/7CzMdUjCrL
xLbdpaVSHdcmKUNPwacxJP03w5H7ZUThY6k4v9nmTCJEr1O4L4hk8ymzdV2d5SX/
uyRy03or7KV9/63l/8/Zv6CvmyXbjmWAVUpsXk/49h3pLs5oZZbvnNaOq2StZ+ux
iKKTk3Zgj5r9NDEM44Y57KfMY0toWP6DZuNUuJ4wzM1Kk0keSRdwFHo9zqOwTrGO
B5GBXPUHMdut1vTdvLY8wm2RE4tv0pMypGrQDFABzjn3Sf+jQesL0VBVJonsUjyd
JO3lKg5OLjt9B8HEdC6f7tqdj36NHo0kSbWwMwOS/2Y4OKgiQFHIXquTkML8AORN
WY5SNbR5UczlBXdYRG4JtjMoAPSntRJwcsWAKwRdtJOx4d5M6iE6V5TQhpBps/a9
ObqFgJ2PqQhCdQ093Qcjbq93RHYoFA6mHH9qUGaQOqMin+z+xymDmeGw4+2L8/FR
abXF5ztZ6hGmrfGyLm6uUmY8NaGRLMR/7FMtfJX/SSFkvLiBNtdGhtjTLy/JodaK
xS0lVW1JpIPAmmU2uO1cmmuHSRf2E7EB/r52N3JbaOj8/sQJFig6kbeX/c4e/apx
fie8E0nV1RBI2TJwqOmUfu9IjPufk0GQNBp3Hm360Xm/ZO5L4WKG/cD4agNY46Mx
V7Z5Z14QrHhuDwGGLnfjhGs1SXLWk6m7Fyld7Bq3BzeCY+tKu3eDk6H0JLyMcQ/P
ChRm/nyuqn5TxMyiJAAD6WRwsuAsZDWEQt46f0CXfdu+Dg4nq93w6xGhQGFuSPiy
K9hgEGvflntoAuIak3SbkoJ1bdjhFoCQIfMik25lR4kOAxzRV1HcSgktpf8YjNDY
rjN8G/KgRpI1Vz36WAPsrsTA1Idsbi+vwqpBtmIEM8bhd4XRK6WeR/LzFlbfmNFQ
WcZSZtk6f/gr4O1/+VuHsCPa098xEREt4v6xrT6cYI5+uxe6guxVfos4swuK0c9c
2pjdl6w4TQkR+LUslBzWSmuQQyMDKfEjVH/ToVaoR1q+1AIWKk49UKvNxZVsLTSP
CFjYyyNCr1qZrcyz0K0KLWBhPFgYUrgqv6H/OjCbCwbwCwYexnboTbaI3pKkXhpc
MdcZID40ctSDkBYrJQBpO1jnysAjuItTSZLX15c62KJeBLL6gNYNQiW68X8pJznF
sh6uRfE1ut4YKPJ/X2H113kI21oX3LoHGoi0kiKPlxtHdD2umgRkyNnaXfbc4iVE
ovG5EnCIUEIJ3ChoUpmz+B6WThDmkUM5/Ljiea0CvCN9sP97aXAksPonW/aW8gVv
S2NaO3MvmCwLYiA0ugFzh0gLL9bhvLovYkeQ9UqdAgdPCvu6XCBM2xXjtJBjggdZ
eB6d7b4s5+UvNzhudLc0asBRTfaeZYpdUt1cUvQBahkqNePmIt+mCFv//PK0L9Jb
6ieLf+toyRrwBZiqkWQ94eZ9BZN9i+jN+ph5ROkWLg6v4pvyQlX9nRveaMluR6tO
WZUe3weu3Rs/X38WXo9WdZfnC4QZAu36V0TbDN9efyzkEhfKH4l6rSKsH1IVesq9
TA/z4sGe8ss+uCnltuXjL44mgwVUMHHQR0l/RYEe3BuYABzio1Elvz72vnHFraV0
OlmMQFGRVfpjVNy6CtbCHCOjbpvxiwC138lfLNGbFsD+IccoxqCvtRgxMbAvIDNb
vcH8kHpo3Di66xC8i3qO+8PfReaHRjaLRn8tizzZHkuutHj8S5I/XWrq8NGSKStF
4w3hN6dgnUfYldprzcjgUMgimCe2pT82pbGNmKhgjnyJcOqQlGHJRNQE5w9LL1VB
npqOWIcwt3JOByx0QSWq59KWssTMinrN8TNhQOMnU4A0STPFdhXrmo58ML/XByLx
gMPd5mzxvKp+ptdVcJUzoj7dEnB2NwJ2xvaEUuT4Q5zzPHHgJeQ/bOKBCLD4EXau
yVmkzJYzZS3lmFhsgjMeHHP1yDbYqyu511vafc8YOMJTqwyWZVdrlPUiQJgv+CC8
Qcx3ml8SoDfooQLuE6UVvR0Qam5/bmLpQx6AspLDWLi1j3W/I6qoWoEO9JxQVM3F
11c27glvRLj1dxGxs1wQAU6ioL7lF8R0wbT7xZbsMpn9sNYYvpHgiYBSqKVT6Ar7
MUm6lTxdio9G9ca8K04L+SxZw/hSkw3s7Gsq5I5x5eYx+X935e0r6lZ9g/oGV+pv
qA/NeiTPuzOLouJ8gRK1m7yjNU9jqbofBNWytRz2FLDkyJHCKdQxuV+chx7G2KJu
05AeFuEwTwMaxQUYQQltjOnymPRoOxT++Ef8PMrbLYTkPf1EfVTEMPcxubQEchAt
3JG85qE0oSRSKZ3xreZyHv2BYkXHPRDyIvpCxdiQ8WkJcJIfuEPurnn9I9EIaiIU
MU5hHmuri6yU2x2zHLafvq31T/nmSuMLoe1ebvtbptsZzMXMd4dUj5hW9eqRWyZw
bITWa8qXhKF+rzIcJjTlMlQdXWdcVCJ5bha+H5tb/tjw6udD3F09MeXwkRQOFHVx
opvOjvNURDLQKyLL0cYP8ZsPB7TYNGlSGMlbzOqZHSCpjR5GMYnM7pep51eS/MRx
7WpRd65rWcu2+Pz78QOme7mWwP2JUOUBIX4rdfT6/pVCaptf1xa4HV3NOy5J3FJZ
pXMWrSH6D05DkGlbWYMzJ4JLOOqsOILzb/MZhsIZPykp3Stch2sILwyqrvNQuQF/
u9BeMRqvHj3C1WLkZ3OhYJg439qcmkrwOfENLeYCOYOaemPsUHnKqPutvit5yYG5
gOH9Ju5bIJZRkeQZUtqX4ayu40dZtm/N//oouaBakPaQL/AKgvGYP2KvVhTGcHft
pgy8L2+L3xor5WSzjzwMU4/1bQDUTyLb0mILPgCJfpwnlnZzVloqgY0MQqQ4L2WS
3BVcDRBKjNSyPcVnlGgCDgO2uB3vV4639jlzk7JnwnQxjwGSaC/r3Hwpe0Uc6pAC
J7qHPp84JtwhFWdO+pnwrMe4c9R9fzGlUrCUk16MOMxIYmnkPJDBIBEQfl9TcGJx
jdFpjNhmAGVoup1ttZFpZD/p5u38A5+QA4uzyklFvBN33UPhTV1yGONbaS21daXZ
TCJDEdDl1E7i+0f4jrr/Ed6jbFCO3p+MzRxxT71khn3TsdC1HEHoDfTGxcoGHDQY
cooH8elLktDJLlMqMXgXr6Rm+mxlDBkmM1nltUZBqkCHwIUZfwankJjDAEGUMjXv

//pragma protect end_data_block
//pragma protect digest_block
HPVrsrLW1kcKS805ChCVVLiIR7Y=
//pragma protect end_digest_block
//pragma protect end_protected
