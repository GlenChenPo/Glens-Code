//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nb3qTroFd7Jprs//sVmCU6IzuZ+OB2VSWa/OpJznoPBxOBpzRIHPeT5WNqt1kxMP
YrCXHzyawnYzzgMvNkS4WUAaazvdekqh1BUgKtLyTsAyWB+AiZRhDW+xMLLsQGK8
TcU1bDlaNeEQQZjluaM1iUOalJNml/b9GJl8JlWytGX0LT/cbl6n5g==
//pragma protect end_key_block
//pragma protect digest_block
uDrVkhScx7ynJOMHvRyvg6dxb9k=
//pragma protect end_digest_block
//pragma protect data_block
ettAsz3Qc14BdnPKT8NHfksWJE02QZEvqRHicAoyk+akcq0YjZq5mnnRoD59s3mO
9kOwa3fBuJI3TEoYDDXVI/SXNYkQVdC41W7clt5TX5pQx+BTOlYfoWdlPVuEtRHO
FYcDFLngX2ZSN9mnvd4qCWr5vezKElZnqg9CF/DCkcxokXU3JEZsCDaYZ7bEJN90
JegBXgSQytZQq6xTBfP2nALc6o50s/Y6Z7aWmGU/+bkYjrjSn8tEcb0j3LriaG08
ToCnB8ReabMND/Nv9s49ri1jP0gnqm4KzuSJ8gX9e71xpQhoHlOkIt8lx2g7Qx6A
jtu1kVOTI0en6b5MXhBlyQ==
//pragma protect end_data_block
//pragma protect digest_block
QCyeAVAMPtkFTsZT4aJvaXUWVs0=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
JOTdfTb8XWAWazitmu+75fOD9y9QjZIXekLLMmbDQMNrdHvzcufrLILSoCHqkxdr
CHiR/qbIaoWqhp4Z/hFmhVQa7i/ZkOPQEcX6bmp2JGGhWrKGWO7vd6xW5tfSKL7G
BfWCMu+YKeQ+Y8J+zJ9HLL32bIw4gVwKGN9q9aGyQwRWdAz9IbvyIQ==
//pragma protect end_key_block
//pragma protect digest_block
y9M+lkNk6f8ri0y+H78NbTYSd74=
//pragma protect end_digest_block
//pragma protect data_block
jEo4kHZWqOnOHoh/4fMhRkZ2wCVccS1jSwgvwAcwNGqMX6gsBDdjrrFYcBaSmw32
Uz2AM/tJrMHWYaMA4wtLRcflPLfVSHB3vdnnhx0QzTFNd9r9JuBRX55CN5iJsV1C
MrtLxDY9+B6zqxJbv/QDvK0keJZlnTQa0GsC0uGBKO/31H3jh7G/5Vd8MY83Ey1J
RJCiiZlrtuQT3pZNwwXWIaLHrKU7Dy2j2CuV7NxrM302F2xfSnnI2CZU357BsqJc
KocKar6aoqP8xK7hK6uz99dqV87jnWUOt0msti9riBrmxd454gtyRYJNLiiTkHiQ
P7QOwOamdvuOBRDbaOyQFg==
//pragma protect end_data_block
//pragma protect digest_block
3/FfqQ8+rh9mR+wqr9TO9w33Ahs=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
g6ZunZYZQCEISatEOHWV2eGiP5dGvYexfGWO3v470oQB9vb9ObZl9JUGAfFNDF6m
QzG/7sGyxSDm6+u5QitEgAgctPeECEtwfG1GizD5Z7d0vqF5FYpA2cJ0bqyN1cYL
MYrYgXDVkmeMH+aapP2/61sY0/6B/nHKp4pDcKoi0mtJhKmvYIl/qQ==
//pragma protect end_key_block
//pragma protect digest_block
SC4sV+NWnwB/J28HvVgxvdFHG8M=
//pragma protect end_digest_block
//pragma protect data_block
TTz8ELmuRxRdqj+9+F+biT6yqB4gPyl8HExI9MWWmnMxcoy8NTn8JPWV0o5LaKLG
e1/mt+OsTxiED9ZVc8BLqpeMSmIMF3UFnHZ3mIWrnT7pY+bPKtiGd42HWmlIfBtu
Yx66XOCZa1pAdNX4j5ATOXyx2RLEXswHyjb2omP8dRC0b3gbUGtuPHPxfwepiYl6
JQ41T5oHOxdaRJkImUtp/iScJw+bCVR16bpLGARd4kg7f1OowyYDRUnstOxYiVQZ
U4rpsn3SjiRiCX62ZvaEr0l1cX80jW1LYlE6xa1cr6SX87dEg9ZOLkHeDEfT8Aqk
J4TqjbkmaexYB8jxn2zSlFi3k0vb4rygpgSGm0ucDNzgUaSQcJ8ZS4IKOhsd2Y+3
UmrqbTbIP1jGKyfI7KuvlVQTl3Jhgs4uM4J18W0UI28mgpSE4vQMgF4zP5n9HJon
e6DzXlpt5zMeN4XidVtYdmUSp595MjibvMMBvbyUFA1NsO4Qklz/LWk52cOX8lt8
Cu/H7z9iqw5iUjXJFgoARtQP74hYhlg5y4B9h4A1ok2OU9uUQ6KqGaP6An1uLUkG
XtpUrZlWUu+07UcxJhhDzrTykdjBaE67ATu4vCImsUziMhGV4vsHgDwDZjdgOTbR
lzfqCTunPzT1ESsgZOYxyAlM0bTWSxnKZuPNzLJvMp7CkCox6YyDBzxjXYgjs2mN
qXo0+xF43uHTg8ir/vs4GCAw3PSG7Tz/bHIknkGOkgQsepieYb1H393te6SW7tmT
55zJ63AMQIs257cc2gqc8+nVP8Ec1sM2ovPghkL6yIMAw23KpONmEjbIkB7/dr7A
2DQe0C5ZSJ3cerbsbju8zwTw4XvxV3h34mtOEse89T8B6FEjR91yMBflI3V9IMHp
vR6tCgz+h3LKceu1BnuBfPJt3XzRU9Tq0FhrSmGgXlm1zZK9L0MoDBkOT41LMG/d
/dlNdh8MfJ3y4TMsGGhkx9TjFOh2rxGGOyXH4eG1MYW4NPjSD4ge5eefV30WwS3z
psVpjDFuBZS0paECNw5U2TETSjUkPQQ7QHUvZaAo/KH3ogXzzzd5D2gRlJYZB9Dm
QenfewAqct2zfEPZDEPT3uR/eBihBwM7oqU3IINfCR3ilFJYJOK2S6fOPvtrIBJh
7NxXLX6Q/ARjJyTe0ep1esgyqL/R/eqhGLiiOvELBDcvB+k3oWYMa+hkQI7ohoD3
cE7tQ/m1oP1v0qGrwEkVLVUy+OopV3a1Xqoa/H5GpiZHgp+bpmrLGHVnM1pDLNPN
4jUq66nzJ3kYV0LWH6QWPkEPUIGVNDofttvhAh49gMBjiwJ3Ipucnzc8VdFFiiKV
EjaXEJ00bG2NgBsTYrJhe7zPBOWb0y5niOBEp9KpeGC23NanBKIFdy20RhWxI+8G
fTSYbLvh6W0XUX/SWXc0GfXiiKl8mK/Yv3Z7npPAF+OOEH28cKNzwBQZKdOmkNWJ
4LywYTp+J3Ds1xGiy0rk1Hm4UReKTXr7XZbovo7QbEsifh/K9QybcUnJubyej1mN
rVQ4UbeWLmKbx/LZxl2e6OtLUwy0D7iphXmrDd907nXj/3lE2LyKa5j+soBYgV+u
Mj/sk/ddK/GT0I3M7X9OyAs/d7opmcHhNQ3YlngRJ2LXGs9tCz7UIAbcPizE6s3V
VQ6uaUZv+AKNwnN+ts3JLucgrAs6ATBSize6c7IqBgUXsEBIejjg/7NeLygEbJgr
eZ0M2utiLVat9Mgmy6Ad/k3RuwOYpcCHBUtTUiJdGmqw4EDhOZsOkGdpgVdb+Hfi
exERXlA0kRStfmPJr+q1i4G60/XgIW7NKO0Vtu54FCT9gqcTJYOcpBJ5wyJ0NipB
ikAOsWHa3iDcmE2O3ZYe3VM9SeH2eNMyk7Y6UWYxibrK2Tgp6OQWX0hlTLV6qDzb
PvKrUk2RnmPjZ3fXK3/OOUtejZmYzBPeRmsDh6FAdRCACXqzQKVUxHRTcq67xvpW
4qLtf0d7SokUTefqG9qK2yvz6Y8mP2DtLY/0iY+Vic1zi6MquPsdOA9+fNtvX1n3
rXPu5TqjSx9gi3so8RVLkuft8oaV1jPnVzrQMwNu8uFTn+kGphnErBORL2ILNDLz
WVQ0naewmoFUr2YslH/L6LkxWDgFvQdlfDZNRgOx2NWY3zIhYduwEgT+KeKD+BBE
bXe2pNfm1omNIccOZa+c2+AgJhx1aCxedjtZpMrVJOqAtTfNUHJVCU97ZjoAdUGv
5lVyqaEt3ZxF4DTaBXxSlqYTPYQPFGNIwOlaeCXWupJiMRiEXzKYRYEOKbRy+jfe
KjzM+5NJfo9vw8A/7h7uEVaD2NpZD/5atwjzDa1TqkELKNPNJgGmB6AXuu9Ef+R4
lV6iR7gv6AKPE8033X48idJO6VbZHNY0OBSJpgn6z/xo0cs9wPvicVv0jwfx1Dn+
NMt6zeyI+S4oaPgSAYjwEozjFVkTmlsfQ1CboqGg5XRk20oXLzEZU+qhsvRgFQKO
bIS5bV1xEO1wH8vl+pplv6vt6emRFMSmzuwj+Voc60eGDjKEHdKNGV/S0p7EH1xw
eMNv0TzW036iexWJycDS3HSB7ZVqOfc0qeCO6HwMyhFme3LEu7kVHKgPlA5yzYz7
chhrUKbTuhvmxRBBwfjF7qPtqtXa5zEGhhVrkv8hgOtAd1Da9LdENfQXvnEuLqyw
Gw01jh9p3OQq0bGWGefPBqG/q2tRK01vG7aWoivQmi+mop4/RXUtFzBqwvlK7Y+X
KM+RoxGnH7FYu9kd9xUOBwtL6hZOHM2x6rBEC3hMDDokv1Efd6h6yRD1FNTS2V5p
vbSsPU418mbD7y4bcDKcpXC4qNHthWrDDwp+TTNx9rzLY1iT0xFk25nTH+PQwDCY
P1LYHxrvBdVDhnNq1aL6FpbpvJxYReOHEf6awzy52/uuYt7ErkJBHN6ctZlYEt0G
XzLQI/f0hWVkfppQfacxmsF7M5QHKJwWxHaP+HtTuaE84eZMSZ69uXiA3OCktvdf
Qg6EQ+n17t0Z+j63JbJwsuHjTbz/QvKb0Ast48F8Z0vov7KDYmHaHko7c+jsQCAh
QOGzE3E7ksDDKfj4cxNSnmuhEkYz+uPXfX2XmE3dbV+6T6/G+wkb1DxCC0rSUuHw
eH++cAK1cUROqtrZ3xxCps/Ls3npq+A6CmUDVKYUHZZNNFbEVX3qwUPSXWp113f2
Pzpa+ptfUkwAp4UmPMsr+IDfNtqC4csXXlFhm1Eb5k5uOFk/YQh0PCEExrLIYnKZ
aGtRvsKgEo/u22UFhIZqEdFMvQQOAWnI2vVw3Y0MTmvPb0ppq34RXCEQ1a5HgXF7
0JSqmtgkH+9DWh5t9/0r0CAmglCWGYeQYYkjzBC9CfN5p6YuK7KR4f62Df+gkRzi
fUwohYLFdvHjUHPB1vRHp174x5bkFhuWHgLgFz0P1ygTCfHZielJQNGKFld3x1fB
RhX1fcOUKozjpF78/E57Uls+Kpc6R2SEzcRs/a2CsD/SwCtvVBrbgrPecfbprqgc
T1oCSpqLdDMEZrAPgsw3r+pIRupATLZM7vZ+ae3LO3c8b9yVPYc7iy0LvRaJblnz
/5+uJa0/7VBmWpLEnnPGecOb7lqdPeNLoCTybH1f5UwJs4rxy6O+A1gG6mct863r
e/Yb3azIReFypfe/szefoJHttjomjIy7jTqUszlt4zZVJjYzagfdWso3iQgFeCfD
lyGrOoA7bm8MOo9+dVqL5vQHtbc8cqwyatYOm4DCfMmZ3EUDP8DxBdSU5W511w7W
C6E99UGIIXenU5qzWH9O4exGYt3TNolQ04u64FxzqqJxmDv+0nnoJPgjcSyrLt10
tcNJMjQF4+Qqh97WaslPUp3CHsKUH+7yTKWX3zJwXlcyNqA/SW/bsTYPtFTnb+33
SQrx7cCrvPfhAYYc6lFh7+oGF/8L0Bgh2WUzMjooHn7QGC5ymfjv5heI/qlydcGY
2Ghf7b0uGA383FzP601lC0g4F5GSNmAm53n0rTOVMQtqXGHNEIsdo6S7WZmzeq68
DSej3Atza9ZzG0HKXakwESo+9xZIgTP3MPJg8oc2aDwmrrRWPXWKR2ec8oyuz/Ha
rjL7ZqbHohjxYJRhKkwxd2fytCZv39aqLpBFxGvVqVrnPHhK6EZVioEcYX72ODh8
T0gMUV+6fJOpE7akHnNMblAwFhMR6D0GVT2S6hrQmc2CZrlDEep65hhsEJ/F6i6W
kibwgt6Ap9Wy9OSDX9yeeMelqsxa2/UHKAt0LDrIGk0OCVucQJWZNE2vwnoJqJoq
4zcZTLj1hKG29xzCOInmbSl6YQ0tG4jHAX+IOxSk+SzR3XDYflR6lYHOxeUZvO9E
agGmnbJ8NcTiFmqcEzAfwve5Ff16bimUiwnIVyF+lL3CMTGWqrtGg+jjYp/BL0d8
aFWIxX2HPsbuuW8oxmAYatX1l3b5pGYWYzYPEJ4pDNZZO+RDhUONb0VBS8XKsUSP
H2gZ6dUn/uewaVUqGx6kPEp6KoWrf49VbCI9U1bxABQ0bx7AL03o/ErR87Rv5wiT
4+OpMxiatmIurhp/6DTbIdYWExgbgh3X4RgUsm1tJxIMfNFKh/GlXnE+2HubzjDL
OnfO3+NdRp5timgGqSTsnsxaRHKChv2AZz+5+ZzK73KZJrExqa5td7PlpLmjVbuj
Jbdf2ehLUwvu7eLaNV+c5WGwk5BNtQ86HelbGmtoIdOVpJV/kR65zsOQuxNWJxhL
ha+1hxxJMzPMivy6zpw+9vpcXSxMhCA4+zgFNBsK/7ewSesKsrgVtvA46P0f/Ia9
cupIeSBoegLr2qGib/P3DZbMwt5fL90hj+4xVi4nkcli5s8c7V/UMR6JvKnjuvHV
3Hq2gTvYe07c6qj7JPnTMnIw9CCVdAvgSPIOzd3EEbLxsrmEK/z3AnOql8zFd5IK
LOfWi9YzdJP6PDFiy7L3dvSdEvNchnKRXbx/Zx1pOmKrhJYUZVF5O/nA8YBFLdmT
uPSftguX/1cXpmXTdkuK4UxbG/knj30m+uc16ue24W169QD9SE1PyrU6nkGwJCc4
Lobpv2B3R4UnZIL1iNYn9K1DQAm5W1tVruvaCB9v464Z/syn25vWRia87QGridL8
PmsnHODKlNGEb+xrh4z26EBaZhrnNpsq2cUPllKNPC7NwnF/czaMNDemFb/mvJG9
65a0Op6/6dsTKf+v77DO9yf7avcja5U5uWKecaIfhiR64mNa8vOdACC7qXDFvRTq
cvnqB1RV+KHsWhY55VjgV3pT02lsE0PHOuF80LdbwE3WRjG+JdyR89ad2NFeFTke
5P9nVVJO32ngDHELAskfILbxo6IndL/XyTMYQtMVmr/Jx66JZ1qm0rv+LlKrijQ5
Ay9IvXvgWKm0FmX1B4NB3d7RfLW9l0n2Fr81b+qggWydT889AWNVkgq1MZ43KLnz
9umnh5tUKWWItcW/9pqm26peSr+/X2IoQ9zzCX0+7ILKPeY7DztuJiefKXhmoZt7
6RV2d8yz5MD2ntiTiXA3S1WRXPAMpsUOAHXhA8JZQxbEytLFZrn8sS5nlfCrq4n6
nC+IGELNjRn3so6KPD4goTL8oNp6RIT9eGk+N23WWVXoWYwCHuuEc2Y0pBluQn5p
njK8R9n+J6b0gzc99b38+lQJ2CqUnvAi1lZZa6uYeQS8LiK0voh5yfqIxcm8j1E0
WgXZ0a42MiPGIpA0S1uWtq0PIOBtSshC1yY/vJLEEr0toe/u7stIhsMebQcR6+z3
sFm8mCtlbOWlWxWG/IAZGKh6xRv1F0CSdU6cz2d7DjmhakZiWZX6YL5YESDLXEhc
N43vp8cV3ZXUV/R5cep+70AeedlnS6nEYU0LpRMluwGEGJjML1hRK3okItrvxI5N
gNhemXEKwdfZ4e9cjWKcTHG7R0Zrv/jvCAKhPRJ80SRcs0N6ZdAAgoI3/DEb3paU
nbo/1f5aKt6Ps/4FeQMPar1XVFfRx/g/iptG/WMoONV8qcXj/31l2yhhXNEHSjSG
lDX1K/wMiZw6dW5kjmwxmlVIuzzcg4rCb6yP8ZFXBYIZTcvJKXyYwMdD0Yyzr+cd
+bmULl/u/6u8OZaoueqZDc4/Z6bLvRzXSsuxk2S7+6IDHjFUCRmYGonVzII3Ozpd
ySZ4ReDdcA9ZmhJdil7HdwEb2Gt286l2z6FVJfRXA09bjxClty11eWgyxRPhHpzz
yMHSpk/6U0DTiS+41M8SgZ8TvwM7VcMOAvm7Z33HrP8O63GplrPXFfHRcFZcBISz
YYTSCqLTc4y8n+hpTAjLxz1qKvPgiw36XhHFS7a4HfQ2rmacFRCHFRxltoHTpK9j
FcGVZXJMAQeqHPeEfgB8UFjGLlObfz7sCce9c3qzDc1lX6Qmq+si8dNAjhj9HUWq
zC1FmjE9CrTi7xwQFb197v23nVZp0NJrZuUigTBSdruERX+LI/4ECQplb+eaoYBB
9xEWZcJ296QZ1g23vNIMkfS1tbMMT8C69ZgqkavzqsgZaexm2N3aeJHmam8r+UB3
EwGNAb+BlMNGFP0MGnY8s+Xc49zOCX1hjCNgT7gSkWldUT51vOoROlmBup2CKT8S
WHQQsjRHtQbLdtjXWU7LezaUgLSHYl+yG0EEO37vXqgSjdTW05XNd4HeOanegMnF
YwyFP2lESvPFSv6QxI1scK7Hd6qU6O3AACGRxnWaX7ArNwJ9W/0Q0gmq945HFieV
dVgzqqdnCcLbTsFQnY2aDK6cmieLLFUcyyqKsvgCtF8wXeJ0l+3f9jPtspNAAklD
oViA2Cp+jGwdwMPb8YpSVXdvyeJ6rAT90mcal3UAgiPEe3iu7SceLhlNpD3eFUV9
hvAigusDbWNCBtPQAz4E2mxC7rT7Bex8Gme1MKJCfQvWGzWU5IuNu33/FmzRL+e5
wT9gpQ9PZmyIqg6c9fFvb8/0KTnwNCPyBW238A1SWsHnRkH/0VnhnRm/UqiZEHfI
RPkaxnigxSVBNJa771cOY31xesEzHDHDq0Ig6oaH0tpqogDRE4mKa8P0UB1hgebG
xNm3w4za/MB8q9KI5YgRfxDwl1lJ/9I3oCXgPSc9ENloskzWbtbzvjTt0cEKGG2a
ElpDa20YKmUNGZV13ddZ/47hA/W6dAd6Rjp5RmEm51x28Wf6M3xfGqSzk0PpoiPB
5vi5TSGiLQC49FLiHWpRUHZ6cdPESzUXBQ2fMmjTvZCG69sN1jc7OA5iz8dACxir
ZTgx2wDhhtGyUz0k987x+WQZh1UWEE0h7Lz+fypxzRt3GvzB8hTq9ci7TJ0doE17
QrxeF8pzldUh6U9bf+mpFHaVa4w/dzIe7NHkidA8cTmJNyw1TUm5cZF0bScQKVRf
C3nbrUDLo8LUmPLlS1SK0v8FF5byb5n3wArz9bK5GQg2iUwghYoXUAKKMMGB3Fu/
+sNEvWdPON1ax7BteZ1P/2lFXfY/fRXB866pmKYK+ZDzP1jhiuThu3lidYDdeoCg
I7WYjF5S5zKi+MlTtcmTRcdTRNFD9k3YGBkjflmAqmmiWFJGgTr0Fi2A1wSQsMGS
r7zRrOY6tVIEUS/sSEducdT7d5vjeaVsdDjqwKMb67pwfMMThTZbk4/opDICBqSl
DxwO1qXHM4yrNjBv/0O/25hGcldLOMLv79WKFbYDQUEIPsgZbxHiK5tinAP1XMpp
eN4c77suq685WmmD5GTUxYVyDB1BOf/0n/o4uYP0Ne5akJI0v5SpqaUdv+T704vZ
7krXAPZLWTBNdAE7V07fq5Rei3F1nQFybNKvV/nfkI5xvj83Cssavrxsnfj+6JSv
nJiMvtHE82hmpk7tv1p04CWuHn7B4QZSmBnvjOea7vJtcYGX5GE4jGdLHknTZgHT
HkuPO9jyUD3O5UNo5fgkcMs1UX5JOVkWGO7VpmZLaDOvn3vl88WEmFvYIM4/s6p7
RqkJ7pdHHKLREVWPXKnEpyaBvjYTylMFUqE9jXW52T80BPLq6CQdHvW3LvigKlCb
rTQKZUhSqq7OiYXYrOHGS3jzfR9RM77w0BLJdSrBZJcl1koY8JccyZ+R8jze8zSY
et3wZhh9tvup10g1lpUt9J4a/0JwVIC6j3faaYSSWSTxrY5PSGYEWxSVHHE7zC9+
FoQxG+83ce62dGnW7gvyyDt88/3ljnBtXxT3of7zGVeqyPD71ROMmlUAiGSMSQWe
dhE5sUnOycxFZVFkoZWQ1yXiPVR0rrMiTUhb17ZO2FCtxC5nRflMP2JH/KCbUuOk
CwpO1/9eGw+cqPRad+QsYmiPJfT4S1jSk4kPga8IUYU7vA4DhHBsWPhugOXRWwgg
Xmo9zAokdtUNpOOgFGhv2/GgxLxyyXC5O1oH10GGaa9U9IzJT099f+6E4Mfs+Jva
N/52/V8DKOoca+ksxEx0EP+XJS+e0pD8kgfWjOVNjmSHgsDVZCZIVaC1wYOUrD3C
/XDGgcIzEMXeb5Xp+dPQHxYwbem5Cn9WV5x0/+8uRuMu2NM3ELIULc0btLGQrNe+
i09iqtaZn/weS4OiNYzL3LLk6JqDsiwCL6dkZMv0MWCK1XJASCFYbE/4ySWKDrhO
aqlBDU/7iQRcPMFty1WsXzBwMuLV8xm0tir0ICORfTXOWx1T4EZlLh88cbX2emAk
O++fcLZ6rhB5O9tqbLR3S6QQAGcyO0it06MOMMVzVis5ng6U/0N3bpq1hGuRCg95
qCdNj2Ez4B2gu1gQ41uuWRx5s/+fibB95N0GUlU4d9LHH1FinEboiTQEyS2aNWkG
eXkGoO3rfmP8NvEnEBusUb0e8jZWd/K60MCL6ca4NR5QCXlp06gPbTaW33VeTcpI
Aj1dFImN8ENdB83Kgf43wRhc2x8MQwjtBxG0fqmDk527GlQJYlbaFzdZ2Kc/SHHz
cKSrQC1oXOseKh+S55HHb7wkDVKkxShWRoAfvS5tCnrrTgjk5FgvtgNGf3ojq2W5
1OM+D4g/Y4NXhj4CBF2dKImHB5KNF6D5yIzqCZAiJkZAp2mlprcTC35Y00QgmQhV
SuPKwP3UiC2rpvhvVD74LA4S7AOV5yB4YWrnaniSe5HZ7OWodMn6RVN5Y2CF+hnw
i+g6EnfQT+LUcDCavfd8FvrGpnWE7a65f/bdmGW3jsr702sL2HwTQv8fByqUi/0B
tYWUvFCLD4gkjzLqtynxAL2NarKSqZaL7L7I6GWvKq7vQtFQeituLY1wXZXaogYK
fq0EnfYwmo8hKXM6NadCYx/E1W95o1h/UCoTeuKKzG7NNO2XB+l8tCZ7HLQ0BorU
vMg04JrUHx07goruqbvP6Y/uDheTGo5+aT+uVXWC2E7fqXbth6NXe1mULFy9fFub
g+pq/kH2C8f1qgQrE6Wt14oIdmNt4uam7f4RvTUF4NnIyYtMSthTqxUsAiw7sQvZ
OwRD94AX0gqWxj2N5SjwBi4wN8b4jDQ/fewyKIeRj+alkuUY42XlHcN+vo/JFd6m
1C2HIEIJCMiZdb2rySgKOPaE+DYLYR4Ivk8UpXByjSY6AaCdclS8tcta7+CHP0hp
Zxt80p3Sf0/mWvRriJ9oO6GCdsxQIm00AheszX0HKUhsFlLwjbSr3kHDsmu6pBUa
OAX6GqWV6mUfXSMyEH2XyD9qWBnbVkXWcBcHSxqAg6mkWfc0UvrPfbSPLvrHwFVe
veCirYPlxD1OZCLAdGn47qp8uerDGcN6TM46iYA3ZRYmNi1LTQIxL+o3Svk3sCNM
ySGqBcwq+2GcVnvmSaa1MrTQrjsvAwspb3VYqhCVY1nrlopYx4vkwq4h4iv0Gucu
J5CAS6wMRoZNf/yw1oJDXOGbQIjqLfiCaR5ESd+OCH7YO25mHRTbMEhkj0Eoaggn
dmAiVBV4ibKO+jNB0T2kD2jJlLOWzRzlrfXib/2O7wNEtUPUl7ctilRhejDadmG9
li2AJOrDdPok0Ypq0TIHbWdxz3+0vRcT/OylEp7jD9F3zoUQsL4CSCNHe6ZF8Vrk
S4ym952EErARGtdAiHTn8Vhmfr5JnWd9843jWXaKImxWLb9Nj7r53iFbIrTlex/9
ti4zKJJuAlMOc3jQCQ88BF/PS1d1+zIARZmul5l9JVJ6LlePOoQ4FvtXewnEexln
jzYaWDEKW4w8h05kICEDakI+USFbPlfZ0XhO322i2r39WZWsmACqo6qlg5g2bGXH
PIC83coBOVJiSxJLKdEN29wGjZPrLvQqDsWjtMQKw79LkttEZrYhulCNFIVbsdkB
WCAGGHjsfiwGX7G1Xx56I8GKNDFqpyjxhWylrf3hddZKl7coZkQn4YJf1VL6Qgqw
gza/dBzFytb6rvVzJOQlsxdGoitnd9zYdyuW2u2L8dlY4/nbcCWSsYWIhmrGfQ2D
L2eLoa0C3VE/FTF8b5zBpLtFDoBuuIjRCrWg6xJAmIPxqLBcAVv7QTDXY4/NTGf/
4M3SEj0CNlaGF4aczeRenzPgLZadPa5WMGNeBjDziRZ1xsI62skv3H7rkBUqZgIy
R0cT/3AN1HcYe6M65BAHNlU1OnibXjt8jNK/IV8Fz/Eq+E7SobCN2hw7583G3qxf
v5DTrSxJSAemXgwzptQzxxfYYHTN1gb20DbqKe6PS2420nXSmPHzHrT1NrY/VY4+
0L3B9MW8PdfhqGhpc4ga7K29/IhGfBS1Pag38+QdhkHGaziMCdmuQ4Xod+yJW57l
bzdfKzfHT3IDDnSIMZ6+Rtcru0mKqOD7Az93163VqnwPDeT2XZf2Ny9TCxsBlMlK
aYzHc9YpPNlxlcqAUzJ1ii3UwXk9iEGyAVHPOIgD6eULGefF7bVcp8Q1sMQ2LLqp
py3thkHnyig3JLLGiO9/hPsDE8rf1pXCN+BuapffVa7veu7/kaI2ySnTyObelm/e
MwTkOMCzixfVyJ3Dwof0ba+dZmQerqDw7Xm4p64eiRLVfZ6ZMWGxsrPzP2GRfmMC
0o7X0Rer7lm5Ci5U+FU8+zdH5h0lRlRRR7vA51cogP3C2GoOoNBvqn9SVqnbt+El
HiYb1v1uL73/S/gekvFR9RHPxUknbMBHwUaSEoCpmyajDcvJPdUlnCRtcGqW7pMC
l7Dgl2lhU1lCK0Vs4m5al4ARiWalMF3javu5EzaSwZPFHNKiHpcS2UVXH1nachB8
xajfsNIlRAD7mCuYzjvAcLa5KDP0e14kLmaQf5LcsuSIy4qNC/gbzDjveCHkonV4
IdFySRNW81YrcGF8/urI9uSzic+wUZH8myWxDorFZRqArPK0il/iEucVikW4B65f
1PFnVFoRhMqH3/UZonA+R9zlBBQGMhbT2f7lncizchMp8enuLLUf73DhLox3juKQ
RSfkzrFAYUJ27O3BIvjMNQkZbKNdtPHyAuXDDrtkU8g+6LgL63kfrUOjmvoNquJy
5FtFn8yuZ64vTCsrLlGZNHjpUWxTYshkFe4Q8IIdDrygoteBa+6ndACXUFXHbL+L
MwdUV2XcRhyP0a+w3Op5Rax3Xas9jDkun6x35GvwmyaxsYUmK7Ay2nPuGhPjGBcR
XcgSARre3r3ducjzrw2Xkn7GcVlWJPbFPxnfS2t1QdXpoozXlT5+V/z8DvRJbjQq
61YRyvPavyVQeqrKX8JcJ5Nbkp42w3Z+r/Dpkus56ko8uheEn3cBFZ+vjbLxiVaL
QKmbegxZfKICUjlsjEPmf0Lx/Uf3N202CCO5ULuT5KUc5//ZTfEBtszmDRCs9BQZ
tvrf+ebocWordzrX2kPRzl4iM+QyYE79fzkL1HdAHhf4Sxup47TJoCzD8PwmNqaL
HKNmlFgCXnDw/0ogF0zn7PaC6SBGrcRKdOz6T2Tr1mPbtSnUV5SwQYZ2ufYHA/Dx
nAR9I8KA/xfcBrgMm5Tt4j4TkOCihCfuPrN/3aIeimAwY8JmE/tt8CGa27IpUuQa
i9rmX+DupqI0sxf8OR0CJ46NtmuyyG4rks5qOh97lGx/1Oj7rQ9qh0jrGBDrQVR9
4EfhNil9PcZzQFlHnULz7o0uZSJXo9f2eO8CZ/lueVecg5IrRv5p9d5N5pw0mWb0
Gi8ZovQJEd5BYpW8mwPsWLdWpAkBOym2HJ6QjZIG6Ph4xM67eMzXdPwvM2ipxTtY
1penoREUwHPBHE6xBbuu8a14akdaX+1d7cJt08LWkWD5lNZ4Z+jChUf5MA3c+qOd
XUsP/6AjODksExf9v4xswFBPj1n56cQUgZ9FjG0JtOZTsbfR96wxR/Y5mtY12/Yn
/BLPLll6JTLt4Q2WJ7vsuvN0cchUGOGLUMFB1d1EtkJPG6INK1eKJmTSbOYO2NKW
FgLyeaz2V9QSp6+sy+4Ulr//bRjMr7YlWUFnvtlj09X8a7IT/VGeqXU2atPKcv0a
byTcj1Whhftrme3VmCZOee7oeMcpApqtLTYPStyHQPcAA5oSd10ilCzHPLRrG95M
npwMXpCK0zR0YnfCLs5A8Zs+Tbh56BI7qH6f0KCr9a8pJSGZ9W1/ip6hTahMj9GB
5pHf0UyeU31ADLG8ELNvYGaGmR89CiZW0WDXecE47vnF0I/W7C6ekTupw5+hGulj
iAQa5E1dvZiZBS9FQnNLDFwBngUaQAd1I6wxtwKykmJ+zsenRIcpoVfIgSMxZOzg
4682UqW827eAm32icrosEYJCFD9JoJE2/OfMU7l0hzJlz3VI9iQTtPFAyZ8lSO1n
HnVHA42BYMwozkf/EfqW7M8NXkPb8oVvKYdU3QndSZOh9nw2SOhACxgC/gLTVW9z
YFa/seLrvrdekLN9Phsb0iqHItTw5x4AnDj0ziBFYH4Ipg2Xr+y2PEw8pbxl4dWZ
7oi2gKqEC0DQIAd+hl4mvomLIzLj91x4vyS8d5yBg5BDnlvcZkqDGMr+Umy1/t3n
RNq9SqGVMnljsEW7AITEk+YTEZ3PfKV72z1cCzfmIuyFhFNJQVNQWWsYWtDmY4R3
KDohZOcHE5cURdDEKPmtQYGN4RPvjae1z0fHkB7JNszHYqWm3VIFtE8/Ht38IK1/
1DvjSDyECmN7UjOOs+d+/cDMNj3MJdczUxsBrKrenUiS2e3Pd2AIkU73zcFLhujw
jK2VxOA7M7z6qfpdnJF+363e+3RqUcedQrPmc2Y1swwqv2lO904oebWQXB1By1Bx
auBKmzdPeEx7sXR9rnOWGoh/Y2s4NQy4OcVEs/JExEOPzneY02bMRuVvAzHqj4yG
4pylnaBPczmHPahDef8K68JuNl/gvqHTyu4yMCmwKt1JDXtNagMm1e9DWyBC6PsK
rH4JMIgXE/fGbXDVvNYJdZSJ6ecjpXzYIAudjueG37UIAEevtFUkd+/W251yuVTT
GZibMCzE7TpnPfj1WKDExc9kicMGcaEf6OY16cBjy21boYmWBz8uDmTSe+1qafWZ
ptKG815wDBCTFiW5GyJYJrdfJMYOkmUwyFJSt8GaGh5hKOJSGmkzeb/O6BDd+WZb
ycnJYSVk2IomRCNXYJewQ8/EZ8weOKFpLG9a4flMJ77k7mVHYDzl2Ga0oBkzDawy
zG5m1NEtQaTzmJ7DXp9V9rTxBhEH0v+qEGZODAnO/nflzhSLRxKWoDxvpYyVjUH5
rLRK9b3PiDAir6I1m2I0MEyiA0NPVoFV7rl/IwCJnSDOrqZBacgqv3Az3t51cbZ/
kn4vJw7jfvstfaQEOXUW/BVYguq3nRnJkF4KpAX/fk9zQ6INzVquAhnkrLNf/+jQ
Y7m090z4NLEDJhGefszXf4Jh/mEibKJD056FtML1W5MvEzuLudJvKPb+YwFPyDrl
G5RKWHrUuFCfpzWO/A/MJZe1bJ1ucZp9DQQ7IC9GjxYNDhej1Z3x54K7wzBp73Sc
RsD19GOkJaensIfj0sMJGooPdLeJvvpGrzSr+iSk7Ya5i9fTdlGy8dM+SK+LDsQS
BUTPDQsT41lkPuReDWNVT1uux+4TmntuUUGJp8hqmfoROalmJi0XEkDTHxcOvQ5f
f3jxR/vHjjUYSQ/2Og0NF7JEk4FgqIeBuVApcJoOhK+YJbDvgQDwMj5VUBYDQ3aM
hjvUhfIq5H/3oCveOLrvQG/ivvjPFSmJj5ZEpeUkrBUDgNcs+N61TfADZIZKum7y
6J12jJjvkx+K9xTmopHtj6rG+J6Wwz5E+xFMsYF+rBeS6R/F0KljdZx9QmwiIRzZ
V4uTRaj6lOCBbTgI15UCpVzVtqVZxtAASvMFvXQoAmsvNWEyNJN5+MqdCWtO+6j7
aa7ExZUmIBGTaPJ0/VpCmJqJNdhzHwrzBmvmzGQa9yqjBQFH0LXzruaka1jUJ1N0
rzjQ5yPYpJ1K+0AZ69NvkAwTITpNGKWKkRPqEz2KGSP1HcXnV3lN2F3BlVb4Fj8j
llGfLyQ+s6Cfm10UKpEJ5tMp9HhtAtU7P60dU5FGaoeHgOruViQ05/7QkUNa0Dzl
s4opwWI7N0ODNScfqgpcdCTyoedUvhp4xJp5jLr99US1wpD5x7iXaTyzzaZdnsha
BNz1ikfSVJiYr+bIFVrmfv/gFH/TJbn8mqnNFGKDmFnpC59atK+tYDw6h9nHusCw
WW2Tuj4QEZR7DluKJuTUhEVCM/ZjmvXvIQbUzH5OItScCFHHJ6lDbw9kO2bjXVVy
w7SZmngoCuTup639lIQuHfGBy+p8qzm9G7rD7dDcAjvLZrBDIW+uzgnpQUefrihy
WMhOf5ZvS/g2ZaUdQJiQcXSC/Zeri5LZKFRDUbU5l0ns2pFdM0WCYcNRDbJdz0hO
i1jfQuGStk03XoSfiP50AJfTgxDuEEauB/ox+tnpKv0r+izk+67dE50yq9xWECX5
9b8tUbJ53hnOvyZQSdFwBmXSN+oOQIZw3rANRaah+9wmM8v3e+m0q6U9nwhIkhbV
WkiofQH6mi3/wAOyYYYzK34MfyqSxXXR84aG8mGEVnMTVpjDc65CgXv9TctMhHAx
AAfgL22kNIQ9kjLFshehAMBp4O3tEZ08ZTxmQtkOZmk18uc1M6BQ4Xnq7xjFpLiv
ZF7189Qkfa8t41YvktypZGM6d15+rNXC+CEi1SjHiOmUd1XVFip6XrDpqHh66C5N
GaquzSmnC7vYBaUKLrbk9erzAV0t8wIaluVGsxslY0+3LgSFu9ebP0FfA+8zUebL
azcIAl5GxY7Jvg/iHX1nRwA/9DfRzEqYq5vKegF8CVAl8aiC1GwhXwg70Uq0Od/p
lT3dyYshis60qDF4TyUVmOPL1liHNbtOMIIyb1TYdNhp3+xQNSxkh+sfnIT5uiln
SL0ADD6330nfG66YOX5IomXvszxhFqi5aH/UUlOIpFSB3TqvTgWU08xn8Ozc/EIC
LqZNfZqZ6mXiu6U14Zrx2FRetfmqM13n31TUZM8xafcKDdJxA3aplWmf8wtvUqcf
M9BgPM2tRafnhfOmUTyWF0ej2WWyRuPOdJi158/yY2tT4fl4KI56laq3q93ymxFA
VsG4YRF2t9gvemD0dJGut0cLkXH4VGVIfRcVkpWlqZiYDGZuIsTpMdbNwkV9oSL6
xr5+l3Uq4nDB7fJ6afGiAtpQRZI70WGkzh0zdzHaZTBXf24FVqwD1FZvA5rp9bxE
SEYscvtcv1vVxA5mnVhBwt7OcSU+Uzhn5WmwTtVIyUyRvp6+D4N48XkAyUkGjfe7
CJd5Wu8Z8iJZr7gQ6C/JwUM6tr3IylGw07D1bE6kWI+oBXcdJn4gNQddL3SPF2wA
SZAJyYTi1NZIjfLKaVLuCxo0+hoVjTH0DWNZ7Dx/mz9Hvua+dl2xsivRYrJE18wF
wGQODXKalthTEj83fNkD4jMwsQwaBeq80o4oNwpZ+FeEkKLz1nJwkUNX4Z4QoA1a
BCfXglrAQQuPa2V2qXHPwGL7bE3ygkLmO8qapf24xE285R7yxYU7XNSVPhpRaiLk
aOjJX4g2LOjZ0047ulp2I+wfGV3Mj+dc1ZOpmbi5OIbNvigwj0TrN2MGAUr7jjSV
SWp0mkgVRg+4JeKPYJ8InoFSCIva67mT3AcrsoqvPgfQqR4c3jmAHgFQ1Se//PdN
UDBQsuRZg+EgdMxWDeqs/90IUjjkouGYR5n4yEpPhcBDcC0wKEn1ZOcHXcCmsKQc
399lc/dUWM4P+q1qnZ0lkdHzcuKn/APYpwh4VTe8Fmy+ktncg37ZWUYdxahTs5Km
TD5x7qvDF/GicVaBf7ijxxFKbAMQBcBCTrpmUXSulA3jnwrIAJvzUwZ8p8soHQ6I
l/fODZmj8/WaBveSTud1MVzr+8too0uwf2UltzfNcjNbZI+5IdEddXjZ8mYuYro2
ecb7DuHmSh5Tva+Wmxt6eENbXQH1kSxaHrfnEdJnR0iAO8ksj8dwNOqMM637jdMK
hp4Fmfykk8GCADYRy+QXk6DTeiDKiTO8T9JGXRpSGZT9FEOI4vgXx6CYv2F6yKmM
CiIV28dfbgUDXEUVKTXXggfCeCqOkega7K/ClLEiqEXV+7jjNGBOS2EUp7T50ukn
pKa8lYmjchEJR996+aIUr4XVtMCZWTbSTD4rmpF2emYs8SNDBOa0mNA5PzWVpSup
Hb1801TR8G3zITVCQKiiE/XrF06j6NOx76nVSS/8HNjxnMlkck7/v3iA3ZDzEGRm
HN7XXjFjt/PAvvnT6/h0EhcLAKH1tE7II3mJv08nG2ddMqNd4u5eYHmCINCeO6EN
Pyr+THqbYwGfStcEzBu6L0DNLdMykhbNcDkaGTMJc2nIKQe7+ftyD0ItyhXOaewh
uXJs8NhWXTx9avYDlBGQZbJYPy78+5uogoJHxhMLnQk9gajcbm5DZCVNnqF6iy3s
mRkfpmw9EoueMdg35FfliWo0ehQV93Mc4iXsGFippkpxdkMjTQTfDJdrZkEGhBGD
oxrGiQnU7vdZlinuPr1nw/TWYnhWI/wj5KJcf8FTUxRB5zWXIemAe/QugBYUCCNg
d8trjiCerzGiclCoCrFMXBDz0mfRRBscBKa/8P7SY3UsDRoqmYL4eo1AT/2SGNOG
qVAhmBDKNdjwrYrlfOPZeSNAWLZg3mcaV+7IX+p9Z2nJ4L2WSW1AFVYGToFjLl2o
XUR7WqnVOrF2cDKKFT7qF0W7C2wwIh8TRxmrpBmnEFwx4vl6GIkkFiB/0hg6uNg4
+rY6zG2IfCBaMqe+BeS1ly9ezlyggFz4jvOkLz8SeFsimExnwBR6pgRXOL8ghtyy
HIUkEhFbTXgBDFNGG7iiV6FfuJTpijrCvVvxbVWMSJP2BTF+BHaLATfoyl14dppV
1C1pxauKGGq+6kG59fZXvQxPySGtXzDNxIYVSV8f4AtBtbxvmG7lwkVJivkqkSmA
H3JjjnT3bbHjNi9J2SaNEIt4DPPmpAGkslZEwvBM6HEcSCI0zVNzNlqx4HsCbLI2
LPFyrz5skG8EcCIvcm0z+lGLyjdHxztvIm4iVW9P6ZMRNLHw0fldE5p597hR3tKt
GSlS+Iyqsg9cDiVG4AGiVIVbOiMODrtlRK8N7J2QYyJmx9pbOZdWWDoxCFPqFa1f
C0boYGOJeQeenTH/3oRONG7DyvfDVambXvZSH3HrrhINXGAF7mK7w746hHmkjxUu
0usDNc6wpJvvc6BYWetzPHWDetN+7NIy3UcAwB1zTW2fHyDRPqmtgREayjwJMHjZ
XGJkGN5ucN1jMUKMPu89eQXvnAXihnBbk7/8E0F0q6OCAZHHum+IaQzaM+OAPPMO
h9XsuY84a3zXfK47SFzDzJKysaBS2tWbem6b62brOJKV9dE0LQ3zXXqj16w4mU2V
QNEYCxg5HYohDTQWSBn1/0klU8Y3JgNf/IyJIf5r2PYLxQ5Cqbx4yAQUzqx23Pro
XF/9i5zjZ86wBKqz/qogrM+NVNQ7H3n/eAsyftWROjBvqVc9l6V4S/cb2m9+k2Dh
17KeOBhNXerjmzaXM2cp43IqkV0pFNUof6RI7QqkiJCQKUUadE193Hnzfw3E9Jw9
qQH6PBKtnj8KArVx1Tv2brNeDt19Tc/rVKveSKf2BpFNb83Pxk/hK422MeXNzjAk
Mi18v0Mb/6fWLOr34M+nw7bKAl97IRNvT0DGEU2REHasgGercT3LAcC+ataaSIT2
xiZ7TIbMIggXLsOeDnOfwl4gyt9RqAKR2qiI3nHRv/S76VbxvpBuKzg/MOR9f/ue
4d9q7iINoKYR1jFEnDz+klClPh+Uv7HnUMW1XRzTy/lnLRutLBXlHG5fBhtHydNd
O/Uqa5F2YitJnfH2imKt3I+CM+tqH6ZGgbB9disfGUdxjVf8Jc7mTva67nReeqqY
elMTPjbv6neJUzqAFaKGiVlKYYfLVgxq61bbNZRYdp7mthXeRRTH1XLf7hp6mD3L
IOKfwA0AfottwIR+fxyThDuzWbFdEAd4WgXhu9qGmHmwuxLYAYsua9joUJBU+3ly
GcQqvT3lFM7UDOtcXBF0dnaHMMktXkwfracbVNmG7976XUSHGSw5krQ/qq8qW+y4
q7dgyiNJngEdx+PcHwN7xECQeFUBiyLdeP1H+xarEfZ7beOwecD8MNijemZ/rHn3
OgvvcYmOeMPOISBpEdLq0IynI8qu6lajs9LOGEwghVkKXgT3eJ5k8zU/vhjHXTRJ
pCQa7GLfr3OofeGuthhALJ1xJexda5ArYMX+AaiwlqqgHbowTXTL+zK34UU4MdwR
p3UhAD+iQLIaiS2jdP8Tejlkysvwt6vV6+sJp7t02L43r/x5+mYYqLDP/OY9r73A
pps3MAFa6BQX/SVZZ9VfenQI/IBHv11dNQ84dpqekF3WeHJ3nq107R/eU0cyCnQJ
/gwV5glYpR9AL+p91PBhHzbfLVJycUs800BF2H+L+isXs0Jfrlfs1No5C2KJjkfq
c7XqwkVzh12l1Y98z3gPJJor++D/vOOFYdU/fPWykiqCxe7b9JzRMLA2IhxP6T5e
CM0vNbHVbQlktSsynElceMBWgT4flBQHxETci04XlPJ7pYeKMf/cYsq+kmslpg0k
23nQ8TQP6JtEBu5PChpm14U6aCsdixtfQCfkDlBF2BtZ6bURWBRYuqSkMqh8s72p
LdzAj3dAjogfM/CA+0HLnx+TQOuINDDVQFaevNZnYUrZFVG1eIQ1xBc8pFydMiTu
lJm2WeavhSUY6ORIb7Vpvz3Jpj2W7SSt8WSLK3zQAhmtEmQulTfnk0IiKbHNk7Cd
+7CUGHC0cuu/JpjkqodHjH8i/2x903GR2nfQox5O1G8JQtHeLvL0IU+TQoaOkeA/
NSA4LpuZ8UY7R2vT37EGqd1HLIUD0I1pRhbOIvO9o9+jMpUDxouUInOuVbdpkjVE
CXPhtdGpLVCIuftk5PVJO7x16BhYtZBbXcYdZfVXsqvf2rupHkg1M3Q4g0JU9OB/
WHzka5lYnYiocfQIs5Uhxu0W/McElsl5RjRQoiDGZKpzAvYnTHxXEF5E41eEr+6L
KRjKVVqzcmGSqU5v3jJl6neR4Us7MPqHYJnNGAYF8epGXiCP8YbHdFc5hFj1kktm
t8pFM7AX3FQWFyVnbCDbU/ro/hPEyziEw1sTyMI2Z83bOWeyzcDdCrLW/QIegu9t
jCtxRi6oXnGi25QogNd6LKxPpjIyNFsnLf5Hm1Qpk9aiixBArI/vozbxERNwUcbr
+S662mftilOebVfOQJiwP5IUalhCdwCy+g9HC4FsHIPkLn9n2FDnZR8MPFFZ7+z9
uRAi7iZvmDFnM+d0SSRw2P4sWrTsFDlch26pg712OrkEm3rRqefCMMJCwRdc34uK
AUiW6SMo/Wp3dTfuV7Lr098sa6RpT2DmALWF6fiTko0T8JIG8T5fXsQ0xelefduT
LrccMe78ezOjZ6YXCnoL3rdwO+RToy5PCxofZricPzZvVf+HkCpUwCASck7h07EA
neX6oZlyxlRPBBieMMB13MTABmnHKqEtCLdcDdUsnb4FC37x4xGV8fq62FiUeAKZ
kBSNgvbfik3lV+Fy3LOfnqKPWXQ6j511SvBkMiPGu8qK5WU0mRzHft2p8GHSiG6P
Boc4EEhpgC1mShxV60rdheOnJWANGmzfEEMyD3Ijo+9g5/+7A5bvmuklHDNt+oPr
pGM0Ahru5Poe30povXUz632WCO76YbGcnDQuDvjwOXOPV6rfmo2eu+8K/dRwo0Pl
iJ36ZAExDz7EYWuqiSVfWSR24YUC6tKTTWUN00bxH5j6+uX0P6wk6Dj+xBPdpVQU
JUUu2ndEHgZG6E7RN6dW7pwtOhpgDuMEha+aod74XCnudC1fDpv+WotrE4OTzzPB
NUfr2ZWOt25SIBEQAD9jIOQflviiLJRqJRnhzLfeZfyDqx4NfuEftHlaHYxfW4nV
bDznvtU87poYDl334HBHnATE6D8ozQLNYkZYllKPmCmtahAANx5vpdP2e2AEZtvq
dWkZBiAmC2L/JU7HPj/bMtCvcSvguty3ejnW+VNWI67VmMf8E5EXveNV0QtG2uMN
Z0gGLke6+CDlYYQjJxhfugwDw9Yxrkay6gWW4t6Cf0CIyAYCdI0OENEJFgiP6avQ
2yeHsfkzMntck8QIZQ/pchqSMIFahv5F/xBPPJrZsTtYmrYcklvFGbS1dEWp80eL
+Sr3N9RQtkez3a5LUOjdw2AefEzSKlULIFAC+EL55USFnevbsJdr4sPGyEfnrQ+0
+rGE9l9M6AOfyN2gBnozTUCftNkQKBPCy28P2+vQEkAMaoOROv2xpuL+C12jK88S
N4mnQ8U8JWwqgxURm+tWlCMga3QkxCKMwX1iQSQqR0InSQIOuRIsO2qY5TSWNomE
HNRsuqWXYoHgtIrUbY21linDULHB5UDSG4Rndn5fEpG2k3CP53ZAMawHrHPmxGOt
01it1Y/UynjM4Mue8faEsrNgRG8DrLcoS+iIUT4LMFPXRJlruB3273jqVSxL47Jt
Y/iACeGSYpthDV+FY3FdIDwR+uc5ElQO1oizyfr2nQv1XdFnK8IpWCWDMcg/bO6P
TzmPIao9AAyw02rJgihPYD3ID2a9Qlpd4wfUuAHHQ+BXlXHMNq1rCuwfdwd4r+jo
8FJu9Jtu+w+ujWCUde+CjJX7uvqt3GKGuXWss9Iq65GIi3Q0qg9lGGhzB9g25aus
iEdzmz91KhexxD2HYXoTRPoOGIb6Yu45F05TMkU6cnKIWCPodPCoNQp0MrOgO27U
5A+7f6fVTN5NGv7MojBChWM2C0y5mzliz6680GIaWboMb61e/Pqsm/6kW5cbsFAz
k3Zf/F+rQTYhWxPHlIi5Pf0RgG48aey5chuHerUCMgDbVmokHOhksPqQ93WSP9Oc
jKVA+WbwmjEA8NNISJbSKrJyjgnP/PRWNvOdKOVVjyCmGHe6/ahiAOoDqBWfbkDY
b+puJ7SQy3tXULrKg1Wp6TdMzEickguhMnzOf5d1oh80L1mvpBNNfRB2+KPrpyBN
cYr7nQXdvEJ8vXV6JFPk+Yg4DKe+xUQRtEmVYnlAg3U4CdFHiuYgPUTNv6H0bYDL
fIMbRVM7Y7GhC8KhTjxjxfPfoYxUZRbLjb9aIblZ3JYY3SMMD3VwjWGYcPT2xMgi
xDbIvJ4A4+pcy6wRjwHxYum3g81JnKqQqex4Z+WxA811Bt+n/WgzjtOTEvCclLFs
Q1CREkR6xI67niWlpIsZfa5wrsiKtGaipHSc/PNZq+NKgXSDQ30R1B49h5a8J7pl
UR6XMq5trhw6wIo5YAYHcsJkWMwX5QWs1t7h5UR33w5nkVb3eNkS920PRvXEFGKy
fqHuXe296qmd3852afKzHK/3mgGfQa5ox2HW/os+fgzBjoEBKZBD3Vr9eUsYOZ91
2EjxSHkBI6u16qZQlkWoCVqPtd+eK3mFMKbOibmEIxWyD+utuTXxNikT8PzEaWaA
XyPn9Q5RE7PSnAiQ4Of4tNBCmj9dQGgoB8VDTyiildhhoo/mZQqYgOhI8/xwTWNo
4m9sgHZR95gMM18y7oVIzldqY487LyYjZG4puroOy3BRVrZjxpNzx1uCwJD0eDEg
ZbMAfP0FNiPoK3gATXGm+ktZ3G4/+jK1sjzs6uNsGkW++UgcuyXomSN6dT9oux2Z
Lw6yvPrmACcpIFJbzEyGeiZLuHmGx6pwdMRkPV00fUZRkF2jFJyz6J7P06MKjyAS
9v04eKluuyFDLEDYQK8M/BS/Cr8rxXv5vuuT0VRij3MVwsk2OkLv/Rn5GFwEkuMu
VZes/YypI/dvOj0M9weUXnrkrbSIl3SczAgyDJK7av1XjrxVEDD5U3iMhSzkuLwq
t17oYDX91Sur0z1m0f+5UP/ilXLy8W3xyd6kRqv0lywu1brwI6AvM3DR+XhR/3Ko
Cm18aC2VGp0P9eELlFEKfrCKPLmH0sdofV4nJogamlcvRrpAqHjOuEsyfj7JckYI
fTuQY15xYpueySVqe61jAtvlleP+ANFiRVZeN+P3+9NNEFpOc4+YPCqpRaS5Cw5b
ES0kZOXs5c0/we7NAKADjsMfYd0InY3RDqejuCcALAmFfvGseuK/LjMYsBi82oV7
PSzY79YClmjQgP1S3X1y7tZh5iGZADJG8mHf9mfDSxYgffSm0DV3TrA5JoQyK5wO
tVmcBQa7tFMzBBkng7JLQVzHBxTFMj530QZ42TQxA3w2UD48TFor6G9zdmHCQ7jN
P28reKqfUUXS+EgpQQCIcSt31kfEGyNJ5L2HTNq+nivl4SAgFbhgUlZaXN+6VI4Q
UCsjpqNEq2jqMAcuWxJVihwvjS01hlRvXOz+tMInLBbjiFx0iviq/Lh5fjInrsEp
ugBdbKa9zaSG6MtV4B4cXNb6lxnqVF5UlChRNlgq8jO98R0MfZyr/Rju0eAk1bMx
cOg3aQGEIvzMl/ZPNhq+ITbE9UDAS50w81yna/4uW5yT5V3CC6bOnoh0soHowyXp
hRdYcGd6c48MGFLqkkeMVzNyegSjufBGCcvFxB+afk5aIpTYIO+OYbIbvTAFHkqk
Y2P9QayVDEJeuWtR2ua4z1ikirIKwvMFBUu9jb8yBVlvKnRoJPL39jUIA4qXxJLn
SnsG/0YpRdaX9ChY4AWUvu/t7q+Cn3/4sX5O9HNeVVrt6G2FV0ZsaCZbHX+veB2H
m9YfL21MHj+OdkB6SJE9GCVEFH8aKzbk0Etv/CNlYETZwSE+u7uUoGbcThuyXYjt
cMRgb5MP6kr6S+MFNFx0aRqEJGdVSecDzuY9rxO4txBgxtYwLUZ6gh9O1t53oVCM
nmoSRlCcZRZXYVB54mVQLnofxD7RyjmDvnOe6FvCWJsGX5xW8ihR1cS+r1amf8IZ
68xntO0AwSY/Gw7wZ+lhrokTqXhhFUCM6Zss5YTtnhMw30eEsD1tu9P6JZozrdKK
CHyJCesHaPLvCZ51TodU8TSj1hWkDGVZxBRsVUAt/FnKyHj8TASlWOPC6snJvTP6
0fvug9UbZ0pJXdnd3dIrsTSdwYZusZ234h4Fbstt6rNWgL79ZzooOQ2yZ/qP0WCL
KVo6kVXh65wR6cau4scmyoGXwtXS2l1sgaR2ke03sNhRs5U0NdIkYiUzyPZhLo8O
mGPfQPFDix4rkz/9r0vkoAu/tfVQ+gWFTBlOEUNeFXgR5UdaHEkvx755vcHQnQqJ
UR+TAwOVsqPdwUedxeTULUKMda10p4gaU4F70+CYmYN36o+XFrm2ASe5e1ifUsfw
gpPfsWHXOljyDCVejUjRZqu4nVczGPxDVBNN9oQWjAW/7aQ1mqFi/gikLYK6l3VX
AgxHCRBDOFm3AGKzP4Elio74u+P0xfCWAASgZuFip1R9lkPW4CrbE2XFTXKGdcOt
GfJIsLaRWdHlq36EIY9k6fXniKy87kYu+SIq8XzTHzFncSvIlWIpeHQ3q2ace/qK
JeZ1rOmz4wgKajS0uyDyqfxyCDTG+lUJ7e3eq8ooam5T0X9RdFwK4HrJXZlLVHcz
kvDI4uM5UwwH1I/trdJQG1mkrYFOwwr0rAC1fXxPmGgPm6J0klo+soVjupPfajCl
bM27ZU0Dks8O6aQhL/oIOV9dld/JRDn2t1M9voRObUw7WQSwj6OElvkPnK8Ic+ln
blrO/MLQshnufA7afCnEYDB2Bsn8NwFC/k3MQDNQaUT/kKQXnEgU5ot7O6y4lfbf
IcnIv/ZaWRXHSbCEMJ2Vu0Uv1xjSMQqRZFeF3WRn34XeVZTMYKsopn5VPNGxhKiP
eEFIS/QKy82vBUJEDh1zb0dJzT/jGekfsxmKWrAp8VKYTuUkN/owCVhfj5qntonw
7tZmKGIXp02YBi21W3fwHhieCARErRgEA8lzQCEqq6LOjdseIGzkjV6fZdJYAmZZ
D8Dppvc7LkzgELywZBRfyVSehMsxA5nHXQSmrRJXjLeCKsH4TKDDxcS2SRJlhwyk
VSA92NwLxwLJAPFR4CIP/YumLqr9lczw8S/1wELEqray7kY23pZaUTcLqKrtYEbJ
lyRwgUOSjLeSgXEgbTQRYDzPZ7Mh15D2jIoepX/LZIFeXo0NtnmfYSFGWjiyqPx9
aXxKxCnJrua+oJqDW9biZkCPTUu5G3kEH52W89tENodMAlkr8KxCbhpeFXVzo2PP
Tq4AnzvK/C22BWs3skZA+uUNZau38dwP3iVAy9IHeEA8jDcdjq6Zzpdh/ht5XZ8J
9tQQbYh2cDzcMOsWilZXYZH2/Vy4zeIpzXDXzekvadC7uaAssGr4KYzP6BcqZTlI
5WO/wdo+WhG9SY9E2G774an9G4Xryb2uCCS7IEDAID5q73vuXtAAbCdgL4ip1O6F
NU6tmL3hbyT4wag8nI5SLBztIWKkcXFV3jIwffaSkU94a0RrrW1aLl3YiIF3ecex
dL865ACAaQ3KsrLJ13xe84fyRs2gaqVndTIBC3B3fv38rTR+bTkUsUI8QwDgdHau
WWUjxgLu8pRaFhV6alj7I1OHtJrQSTmNhdnS2WvxsOprXZtB8QaVDjPjt37ewuPF
Q2yoIwSVtxbm70XLw+cwI+e6EZhUV3wcRsbS4bEuymYbtYks8r8vKYHGH0hcyZkA
2dlf0sEMnIodxZVjp+6rkZJcO4UT8xUgKCzOoB1NpRWn+DWc3ignzBbMoeTOsTbF
MhFyUl3Kl3alJRHjn55YOz9ZATSgQU9LnQ9LeN4zlUkSJrCULtSrEMbygGw1Tmyb
okCAXaFIKinf+IhYh3bPVdq4GJ/KB5wnFFuTZz3o4v5KIQ9B/h27b04vsOFzrRLW
4luZJSbdKwZKItAWMilAUFF9SfJ5nHN8+7tRqARLEwb+lYzi1J3D+Y7FrjtjKiOa
OUeTcD6mwVRlWzulw03kbIRH8fTsZDOOJs7icksT/jmS65vepexpYnYkl3HAc2Fw
UqsFalsjxfSqwBILtLFYOcNWnZ9tZgy23zdDtqRltj6+O3dVYanw5wcaCwX0ZQZk
KQ5RMYztqDZq5Yer6s8/k72AziXGy41cfpiV9ogv/DWRiXsJTgip6MuUmeQfJDlF
8NrvxS0QQWKdEXn4S874inq3TIilIb3xn9hJgbbMjFIPBJA8IrG0XyEB9CHk7Y5v
3Av2ro56VcSSF5rWoIKnj4D8sHxeYAEK2abOerLVedctZ0LTbNFv5cLizsJ14BrR
wm6MtFSxymCNn/j416zDmL140fi4Jl3bcNlrsk8oy3iXuW6SvgZqIaTiabeFQxwK
XDTDDZllLpVULwoINWbXzU9QepcTsZrzA8ef9o40aSMgznywaSR+vfwoTbiQrWNd
zv+z6/ziB8vsGS6/ThfXmDPhzCAQ5LjM/6vhpOgA1hS7xRnIq583yRMiZY9mCWxe
4c5x6yCB85IKfgVBEPh30Ei0LxnKizzECUeo8D/CgcbvT1jrAIC6v+fr7gDr0QAF
p2nTV0t3GGjxVJcpmRyFRbi9zvkCi0EWnQui+QuXA8uqoDkkbnnWKD4Ajj+XBcKu
yoGebO6qG/sJc6JJqzO79pIFs7QKB9eC5EF8v8yZG74x63alhxOtyMdNhkMtpbpH
43cFnCH45R8qbazrBvI6FVC1e118xmrgj4hxT/hp5jkgqIwaTqHGh8x+DBtArLxn
gVsBWnLAAv79gVv2nlqu400TZrFGgYXZZWKxRoFoKSxQQCecq4GvQO6QmaMz/ACl
/4kv4XuR2yLG+Ej+P07yuSTKBtl8QQ+8pDcwCJOVXHu7RodcSbyrkrilgjM7iqkP
PD6f2vfJgKJCNVyduvOGv5RrDD52JRBfo74O+wndEHEUNwZ3p6swjb2oPkEja+49
thFhLGmeadh+xgyl3du51ARTrU/o62FN6K7+/m1pgBrWH/NRpwaRudFMjVULQV28
GX5X9eAvFGZEnjtzstLlTExUnwUsGt8G5h7Q0r7dnMmQuJiVgO/LElzLtuLx3DfJ
MVxB0fYvD52zoWLkXOJrr2dzRqDlPeiagrQiuuU/KldXIVQqm627UEftrJgjcvxy
tsywaBV8oW0tf4UMVpaxC2pa0dKPg5ZWBQYnaVruPa1pUyiLhsJykzaE5Bw96HHn
/vtiVyEyfCLubIpK9cPsmNDG6M9Ice2SMyHhXxWHxquGhtBJ5UVXgW5LGmjo5ksp
2R/amXy1r0OlA85aB5nBxu6Q3O9C9Qk99rHdIHOlFpeA7zddJAnV3D1te8w7cbgz
slz1Y/EWpDRZJgvPV+xFJQK6EsonUOC1jmBoukhJItWoJTU3rKeIThMXZTDVUfiy
7WNHi8OvVr3m0euQlXa+adL9fFz33YJOQqt7VXjzf/OadZ0UGH4j0bGEiBbOAhwV
iFLBP8YUxkPw60tNGoxVzFj8ZLfVjJBtL1GQYoz+z289yljvMah9naN+hVTt9eNa
JQYHWnZVuq1yHq4ZGrwCEmwXLHnHF+5/PLhDnzu22thgWRhhiNs3vH4M9tujbaaL
0FVFj4qSIWm7jQLShc9qZPrh+z/cDQMYiUoyP+qsz7kIBNWgNoBUaS6EJoUAFIb5
3TrerPZE3oXR0WRyznQY0+U1LYamGpOGUGzHNiP6zEfW88g1/XsGN6LSY3h7qLap
lV1nr29W70Hlt6WGbNt0oAnXTwgAqoystYwwyJW8c4bJ47EnKjasCI5EKdvNFEA0
84kNCPQb3szdAEIKAWtfaZl+1v/pVVRzArsXtB9ojg0bf17gN60vCyT72ip8NgyQ
uucd9Wc81X//+Wt23v/ZwT2c6RrZe+M6XtnvfTupZcbV1HdJB7673q+k2AfD5R1u
ofOEwCT54lDtb2RwcYrssVigslBd9Kv7PvkxAaD3Anmq2zimM0em2+M6x8t0AO4H
n5LeJq/gM+cwSbL8QVzz6pa1I5+kA5ataggj+6Cuc/yB3EsBmWO0sRNoAnL89Nyx
uARN5p43PQSXD9dSo1NBhUphw/6SpqnXh/Ux67MgcrdOLjNNLK3XcbYDOR/WYwPM
bvFV2d7sSwV9G0ZUx4HpWt8bHFr/YtT3xHVHYxJpmCvZwbUzjKMAJ1N6jmCCPYPt
q+74ROQ/rh540do4EkPbZOYCkQZ7dqQAjjfnyLsucR/xySfm5ls6sANoV7F5IJ79
NUNmDKYQwPRSqtNGCEIep6s3uXgSWr4NK7B4PX5NzCizq6oAD+jx+S/lsvpXQzwf
+Og3lsRYbXWXX3fcHT/ESmgEY7uohxtNRbVjuakjXFVjqfRje4EEZvTtkwMqy8Px
G12jnNOoyj0jB+8q3a7MAb+3t0dPpUixE9PrHFdzQbuzmudc809OeCbMsOhdBNDp
UDCuJwduDzf3svK7KtF2gQQ0Nzd8cdlB/wjEXk0LbFkCcc3y5LkZ5dFHlvKrlxMQ
9wnRMII6darrcFyBZy1t9TRbXlsYeRe3mBOIHduiuDy02MpR5gRd6sOOyYL3AE61
VauEijqt6GHgNrt+4aEF3xZGtfM4IsoyIvLqu1oC6e/lLxEEpVs2fsB+4jdN3EFF
pjXo5gNFcuzqQqhyaCvosWtpAOnNPWSSrebo9Xo3ZrRgYYC+u6po2xSbSdWknKmU
H+GQNwKPh7rnCLXw10Ee7AM61Uj9bZWN3DWlLUPX+LAcTr0p48uckjEG3LJ1k7nh
K06ivj/CgxV4EmyjBsSWEvucQ/MkP73ofT+WXgTnelbFrukuNwPIbTYuYhTAnjZZ
sD73WIAtMHDcsRTLp0/BvefD83nbBvgyqa1u33gSgE+cCwgZ+FqaM7GiuC+fxYN2
48SKpOQGH1YD7nC/v0irBjhS6cYWwOXGCfFtQ/0U/lY1dqwNr7IHIcf5bnmqR9jx
qJdbo2TP5z5nY7i6/GXQwknE1qBDNCai4ims5OxNcBfYPL2dXFDNHAtYQZrCNF6g
EwDHT8LHKM/SoqL5aMicEsn1V5NP0s4v5qCl+X1DsgSVvwFOvPouxZ2wmTsdzl4n
72t4Jd9pN+J5zu/6rD0B6QM7ZgCRG1JMrw6MbDpsaCTIoGQSivBt7nBGoAkqzTze
xfXtcGnoCb0/y9prLHWB/xWyGbDBQmk5RF47jf6tEbm2ecBMbzNxN8/vd+yzZKNq
0quKRm8COl1Oi4ZNkjDiy5VoC1gEfRMNQ7JfbDZz8x6uiN4/C9l3S4IGG5IO0FJF
xInzUL4Uv+LDb7I/JtcK97cTUwJPb9VWj6eNsiOLD1gGQDrGzw1iBYRKCaW+ort3
aPW45G33eo1AQ3+0Xo1ruhwuTkVWHX5djmcc3MyxkK7wPcACckMkKUlGV98s9HIb
vDHg6ksbxjrOFKv6ZrWkNhN3idakrqrDJqEZQwwAsF7OIVYBN3pcw6hTLECi86Tf
cAdOSX7gFkeMMYmMU3MRuSh7O26tr7TxGpzlxkD9aP9OlHzn750SAYBgKrlI1KsH
4ZTSyPbzQyKcT3IdVKxpH7dapKBZ1bloh/6LmDnruw+eMXTnhqdyqn4omHIYpkED
TV8LOSOV1o5cT3p9XRVPzXCLwYz/kmX/m4X6DOZeyTg+yDIr/pKMXacqP1yBmJ/T
n1tXqJCeWOiEo7sEIJVASGv2tOBAeScQZGEUJ+gg27aprEs48HSXP0AKRxhfWhp0
Q6K6m3vxDnoy/l5ESqKmaSZrxgg7cMzLpDf/9ld1RoDsG3kHm4uU24olZW7vYqIa
xPipaTpne4mSvkAOgQOj0BYdlHW6GfFNUKfskNryfX9b+X1ZZdAzobs1uJl3+dRu
BGAYRTgHHTSPaZPKIueKEtuztaNkV2LjkOgYrJWypyTgROjpaHOyrmdUFB5ga1fW
s5vsFJt89rsqclzelcbUQ1TkhUAZ7eKJlKCefMSXObMI+FkDPoj3h667WTUyc3yc
4nKv7+YbRBb1NvS9H+9PbaXDxNCdp1MWAwzH0BL1XCmCjEl3LIOWwun573efC0n2
j3bCE1Q9IpLmNFjvpCJvivBN5lTQWZJVtEQ/ConeTYz1BWg77baCogh9cFYHs7J+
f1gJVNjESVZ85mfPHuyEeVo/PBHOQ46R036P09foXyByz0gWes5hzJ/vr5wgQo2R
RNj/C7LV2dsHduRZQK5s67WwKcXYrBt0etJtnujPsK36eos5dMhFrY08W3CaqEDJ
weH/pLlOCYbWnesvTQrGCwUDXfcb90S3Wit/GTqd9whngifchJ6fCmokUNofjcXD
1tIuTEvVDWfVQ3kNha+tEcWSDgMmmqAuEsg3yLc62lEPcpVw3BsLVpo7VPFMvi0M
m21/RkOyiGXEp3eMPpJ3nPVUS+SZBUZmXHKau1Y3CBNLOGW3Uw2rJqW8cijwFlSW
G2CxdCdTAeOPEGzbrH+DPYBQvCINYTxqXmE3EsBbI9ykLrBm8elt7nTmVETlS/fb
5i9+w1XEsWQEeScmhKb0z99RsRQ+fRAjOYgQVq1PWaiA6XoKRbJZon5Thh2DjPNj
F0cMHuLWZDpk60G68dshsLwZfvTvQ6EokqhCQknJARTDBXPV8HU8JVUnggI+Fx+i
dzuPhlYbGVj4ifdzHN7zDVGSLoWUFEOIlGh9eP3TBxpI8dqOs8zjgpfvJCCQ+BJI
ddIZkKMDKjIK9Utilufuwj2cX310Y50a9gprP71XTL8n368XDZ4hrUiDmKZrfDPV
POv5fW2CqMJrMyjI3l4A9DaOMGMI0s5dNoLTZnFjU+ocV8XhOEDSDf3aPnPTFTq7
3w35AIycc9aJCjYggofaRPE7fuLODeNXjoz/c6+SukXdA2WAgEc2qsmGJB7cmjk1
DXT/f2v7fYxBmvPJrVQFT+s/N2esN2fwIxNE/0grMZJB33DGDyDgGdRRxfaGjeXB
Nvoqrv5+ln/T1I2DE7BypUv7uVhdZysHFMV92szTYQG6NVxWFtTkr5GDGlglmS8v
/WyyUY9QYNbyxPDELeX7g9CeycpMMW8lgQbFlGREGqCYHidwg8tVvMSF45+8v/e3
7N5h5C7aWHRCkPFXI4lG46uayt2C9JbagR+vffQzSGtCFy+Ep/9VgrkLXF3kiGOo
VEG0tW72OpPe7FUBlnFCD549nISb2/rKtQLXtOuPnoGjQtR79NxrPiHH/GhK1sE9
ICaCTr+IGh+zbcTO0drbYX3GR3m06+sqf8zrTYX3jWah4MQ4s8RnML7mkDEYdikl
7Sv6PnEleyduDYvTFyccpEo5lhgLHBEst4UT6Fk1R6Nt1hwEqKw4Dxl/1VSz8WFs
aHHOuvET2ttkKhgcVQetl3dS+mZc6G8jcgr4/i405sWgZG10SBSi1suOizLqMCyX
Exv3RW02totY3J1SdeQhtjNGqT6CRXmh8sdkqgb0lFrJi4fyWyp3W24wkjzssoOM
jwpWYSkEE4UPSZ/rBr9UoG3Ob3CskRDdfU0QF/ouq8jWVVcF37UphNa78Q1VoMTQ
4YFK6JAGrS71KDzY+b9pD2TC/DWhUZr1KILYg6Hgy4hJQwJmb0dAAxX5DfY/bwWg
2W/s502b7MWHJL277TOLV1kpiGKWgffauP7N2kpyDB9yHdx2SPd9EHROuI1MVfNG
0+9d962Is6uDvb1OUfQrs8DXtB2PtlpNSvmzmiOnZOIC/xkmsMGQXZUgeOIgkLT7
Qr3Dofarvd2FFY3nrLneRa1Q550NrN307iqODnHjekwduooBlrKlVZVhzfrPeOiu
D/ocS4FTp5Q+bvrIPjta56cl4bgz3JUJH+mNbQHtpUU1Ct8u1i4Zop7MafBIyOwS
DCqv6boQmM8l5HeUIJn9GBOmFJaKJH65q0mb9gOri5gdKET/pzoj1Nm9EgHja9X3
lJj/oi7vd6t01zXVXGyVEeEQZvH2sNJPFYYGMgAEvf1XyL+uQbZjLffra62G8oqb
tdLvIGkyspjPMOmAI4jBLuw4ndTABY+GESEuohx+rrnfhQOEmpUTIjGD3saplaH9
V3LCT9QXBOXua1om07SkudC4RX2PPjMl7ckD0xHthptm407Er2g81of7alP/P0pr
KimaZyUd+PMpfNi40Fe/nHJA7G3QHsBBjn/bQTJtVAfrwtNpYaoI8d4uIb+H/7Cb
hiXdMlAZVDUM31Q2AjZS/cktLpN9oSV24mBh3KPDa8OQY4OpL1U5vmUxxsrs/D3e
E2J4Jfgnl30FGRif5lRZRC+U8QHtL9QbhR5qBCKnNI2vkYtjcFL4Y2uBvkqe1HzU
K++aZ0lJT/F3PixpKnC+upWCJjRF5QsUy8S36NEiW1BZdEZwn+xPNJ4IKfoORyXy
7vbSzwuHAKosxBJjUBh4DPjaGtv8Y1fv7YVfylRuAwqyG4UHYun+AvyNS6qTTkWO
CyGl9vVl0K1ZWRaCgmTfdDL4zfIzMFOf40HjGRjD2fnpN/WxDZtxHWns0JbtPecL
hcl9FUL16xlBwRZkR5VKvJn4tooz7ZS0w0zncFbjSLVGaD+vqWewtO/kCceenuZw
g49lqLJjsAlR8ExxRTWhAgb2zsrgS26u4rWuRvhVMxoiF5x7y/nMCa9syU6JUyaV
6XMFLv0YUr+z7c7q1s0hov2eaFvEmuf5ZB7STYiKE6lRgAmJ1mo4ESAcKw2B9Afc
F/zy78984KPRsAyIBTmVGIAkn1sei5fFQNM3N5csXWIxgiM9s+QSM8yMVTPPRxr6
ArEUxCmeY4hj2goI1Oa+vJNimaW78n9oBRmAsC8weJ0xsHNDCvPVGcJygcJGCtV5
kP0il0Poo4S3p2GanmE9/rYJqFenxvEbsyaGD+58kB1fM9dLuv8zEX7M4/iVBdAm
B2pam/vfJEHzAIjw4oG7XGgUnBJEvwDBYvJc52rlP8cg0p0O4Iics4Eq1BMq8NQY
yiFV+WuMLgLpt3ldoEXkjN1tjmaJs2pcpI+2uJTH/izdBwoyZTfNFpizrVPFGPkZ
zqzmIl1+NT941YQKbB4/xskbFb1o7+tWADomr1RmbfmUg8hGdFHrW13NzTAGaqVn
P+dgADhONbXSNz03gw7PnPFjPXmV1qtbBljn6DILYHE6vsjQmHX5mpBa4vWWAyKi
qXdtI6IYxi1kgCu8gbfuX19vjrwFKp2muJk/ayZ+iEZ+9PLlb1dbxfyICdv/6Lax
MaCIoMAc8+N+TEIAgNr44l1/aGJNPPVOlS70EDvKGhDrljAFsaB9RcPdKxFQUBnO
7PP2Nh8QluUVqnHUQwIHUURJFo1+bxyihuH9RQR6YqmCKiG/gULf3JetH/daBHmY
/BttNr/tWm6rajKuH4D3Oy4QYa9Fimpn3PHRkQgKbprRhdGjP4f12Zno7smPFSbp
8VRlseTKNl86/UESpOqOb+4rRhnfQ8O6Yy5f4Ln0qkVxpvvvO3HpooJKHekek0mM
zSfGa5Ozn5r6gjbgBzIHQc5wXfSoHMne4ymNaQ2PBi92bG0YfQ9DtG9/6gPD74WY
dmf6iOQUcdOhggpWRnQarccDTMe9gvbmIY4zEhggK/YW/ue6y2WmoDimTtBFDQdv
pN1N9trjfjHRddJIroWRZzRxYqjF60evQQY6VrgWWQhmT81YudOfcVrFE2vvq0cg
QfSZ8KS9P1HBCt8z3pgWuLv5BphzrHL1tFnAtlxvO32XDLojTQ3YS8gkbJEDoqmQ
1TC3UjbqGdg7Zvx9jfPYsoOe/aROblVPkot7lCEltWFuAdIvGh53akkftZ4pbLZM
+4qJoeE9ruPuoBTQAzUWO//zlvmxg8EWXmzrupdCrblPC/t6zxG9EpjnjEMAEedW
xoIS8DsAsq+u6MUhChuP+EPAU2uIL5uwXTce64mOoV8r2Iznl7WCzFZDA6/YLNgJ
CB5DoxZ/CxA/EVohGDwdS5sehCcQBX1eyBYH+3kbhPjPVwXoSxOPHo3iz85HXmBm
wcHP5XgCiXuNtydfwXOLoRoVqUu8iTb9l7y+ZEeDcnanBW+Be61jyyVWoXcSH4e7
UJ5R6Heb0nUxAjXJP+6+QhzjuWmTRMaJ0+wvAjndMGwFTLQu6QqK+3dJ5M282ZVY
4TgCBCWs5MdZXhXutBejO3p8YRiVLI0WzfKt/vuXRoEecRJlMlbDuFyUIidkXc3z
cRumDLjaiFEYezCngdr7rzlad7uTJq2pfOsGQgaUcGF/J2J63ZYKJPO4mjaQKBjp
oWdWf3g2O+uqy5iAJ19wxSofMU7ZH7tehHJtUoE76EFhGCTrAteUxji2CVnW0PVq
PlO2sWCCzpzpXu0NdOKQBS9f//uO8+bakpHctpOcwn6/s1QeJvWGUyFU1PdTjHpB
92/6pUwFJohNg80XGFLlT9O64lDXQuvc+Ds4LPV3ENI+o6o2uxhCScpMB8tZIx0u
0H+6E4NXr5gAXg9Kt18cT9dQsVTiRQd74AnqlkoyWM53fPE4anj8xue1b40BJdHs
dhplEszmPLjtLjO98QDZKlcxjHPEj3O4v8qH0ydY2YohxGSDriVYLIn67ZHQqvcU
lKsFjpjDNYNPtwpNApWlGnmfsSuKZpSXGp58lu+HJQ1YYjMevMzwN9btO9NuQg6a
oPSla6+qmgX9B7Uupz2+WfpEeqFkrOPARtnrxpQuPjM90wPrSKN1/w4H7VnXnKkF
0eN03pLMlah59i+qpiT7W6bdf6C19yEDF8yMj3V2EFytg4Ry9RuSRq7zRkWhrhEp
/QllsBW7AmdoM1em/CI+xTaI09O6jlECg9AVRGuC+VHA4ExrwPcbfDft/08PKIVj
oKpqKhCwpwQgT133MdwMmSP8LsWu7aJVA5kG57OHFJ6bZLrsL3Hfv4buCNpKPQjq
gpFTIJ7AZugKVu/Qgtc7HSyDqXbqVC7QDLCZ4tEZv2LOErlsE2fuwIEvmfj9A+EN
cLMW1UXMdH6RjF1fagS044u95DAQdNlsjSe+QYRPCxR8RDI7zvDqkunf/WfUJGRC
KXWIRxJQkzl/6woGRiofc1dDdLmOxFsoaNo0WQa22alLwXmzIMy3a9Vr0hk4qgOm
IYSkwQeCH2oEx+XeYqtlnYhKAlMXEMelvWqJ6dSP6h8rk+2RRBSL4DStuxXmUQ9J
i14WaXj0+krMb/QOyftLFg9ZwZcWPUATUDzEj9U8BE2SxqCDPvh/X78G5YDti6YU
sCd4XuBhZ+lrfz3DJdLU1GpEb9OFRxgTyhMDBaknr20uch94FBuBNdNvKckH3TTK
pW8vxw1MNe1V8uFFTqjHO8FdWWqE/GfHxF8XvZ0emH7Tje8IGYVVVrjnoKBy5JLN
03FmjHYEXR5JYk34l4Q4aEvE9JoeBkPuIXfC9NdrPIR4GCWKnzzOoRekI2lVRvnp
iM9DEbMZtjtH5lfTxZVYnTHPNGi/k6JbONteDDqztkNQ4ksv/L+oxwX3x6MHpsHN
nkR0ISySyMHJhUUHIoGrP9JwRqO1a2egsEgLRPdfNb3tKaqLHK148mXrtCTNjSsd
vsJtljW+xziWH67S3lTvTVD4gU/tlPirXg96WN8plg8Ci19Yi3e4k32FIxPIuPro
+PcVSpsh7w94IUBmwSNhfJhUZvJR+5lzDGfOE1NpSNPKxBySl+Ng0jLUL8wzt3bE
5GGJXtCoSZWcVpipa3YPp9wGvNv19H0Vln4hMlzGeFhG/VJLw7rDY5AP3D+T5DM4
r1R7OHpkg9wxDKI1ZVj9LLSnf2OWUqqr7hZ5QM31PP92ajHC6q1ZOWe3rInTePuf
fRh1/05o6xPHk4AK0eAdmlKRSYG4KmyOtnUM7qWPIIEs1UHDI/V2jl7px3XbpVyE
fWh2KbHPCsrVvmM00wNmW183Z16qzm3IZ2bhBujb2OGXYFnSQOskU9DziO4f9jOQ
RFDTu1oBZ8fDURMRU8RqlItDdyr4DwCaMV+om8CcRhVsE0g+MMG54ALgmMQvaEgn
UgXsiJhh8pruZ6jYKeCs2ez6Ke2aNm4/WlRHsnzOTDdiundfGylKDq5FCUgYqDtb
u13K62wUdENOQumjYAF7xY+oY15k786HG1jIs6BEqbyasozETlJy+Jfhw+d9ue9+
ws0WnkVwYkhhZr/BOTFa1SKggu8RhOoDVN9oFYo5nREqUBY94V1SVviKw19MHdi/
43gGJDgZJRs9aeAZDc6tawmRTmjpMOZkkcFN69kVLXfEY6PscYdg1H4xEuJyabFV
9ma7pwH4jTQp59PQRtKTbN3iSZw9T9ySqhnoixfBeXH0RA/dn256f9qVZwMX2bcl
ZtP+2ZtfiCjv18KmxrpgmMQ5/xiclxCekEKlYLGUoDKk1U4NDV7ui0w1VCDNmTaq
u8jCVlCYbx2aRp3SAUbVjOgbD+t6UIpxq//4Uar6U1u56CM59Yx7IWS+iyQp/nZ6
umxq+7hxdVWaqeNuIQ8uUSRlbqhC6fccjPe0vDrGdfBuVnFdaXpPGWb6GNbKkFTp
4sAbHby15NfjQe1WNzoG1UO+P70aIs+hzZ36GOj3mIQ4iLxFMblXOX2zBzQeFM7Q
CEF9xgnTW+JQxulG2U15rFAGf9bWc2y3HzOR4UyJo53f3NDotOVT0PxBPDH++W86
oa25icI00jZp1K9YZUkFF7aCNlqiRqEet8w7TuIZCfo9jgfzbg+fNrZLqBoaLtNA
YFd3y+fyFn0thFT6i8xBJAKtFkFTt5QSMtlVqjJTjXsrcy70K75jgY7Ptk1d1I2M
P79IiEIUQW28k1rQUf4ebMVPpLaxropjFiRm+bqPNdiI2mM10EFoBeyEC/ZkA6Ee
GvGGUIakBddMqrexu4fH2PANfuXFV0Y9tgq8uQb6OMUCbqRMFkISfyIQ+J6glRzt
+h9WEjRANLv0QW8JLpJzj4thPshoT9MGgs78zj3EnBKR3p4cPXxdslogp+dkO4kk
0N0Ja257l0Fok4u03Sh3h6Wz+GZj6arUnsMty9bRGpwUtOzxYMzgJp1ONuuj06ZF
QG0lDA64DPv9gvRn5jLpaqP7yeQp6nXthnvsDZqExofCz6hO9WNeeSEqZt6XiZHK
2iDYnsijOCxKPI1BfZ0poGu2tOXlTN+J6M1rnbbfDsIGGGaTPLa4w51s5cGO6VrW
34INt9ffqQBCaEvvE9UI8niaqNNRP7CfRHoY+bzsQFUG1ka7eEmAnnp+17YxlTi7
D7FSOCTtsrGMz7jbvbl923I+LMgdYg7jyRhurG3k1az6B7ZTLMBIn2yknxqMAruq
R7vwlDKmZoUgrv+dpTqB+ALObG8UYQDUwU1XHCmQzFPgXB9KU8qRelACTEL/DA59
tCmJPyrvoqj3EABLIk+AzFWb0lv/f8i6/eJSEp/aG1+oZuixDecDk0o7AVXOdXcE
6RKGbHTTbZmVnLRGALzz2v+ldbgkNM1XofhYkg70o/G6DRgZ/56cW9gjS8a1JGxQ
u0eJpuw57wfMBYwZwa62w6NL7hz+2mBbijkGCiSGBuROzKK50twD/xh46Tt1sV8t
QeZ+QrvK/3VQzlji1nXsoujutmvVUXXEoUC7CZgL+CThvsVSjfYJLQx3vj1IysGu
T92DLEO11osqcRd2Dssstv/M8tN/A/YF7jnnHrO2DLjqodyQHHK/5kgguEhAg+Vu
8lX/n/8FwKsUJLh/erH0KJRhuxLjAZ4M6KeyMoxwSLlG1RwgUlQBnuZOmGjoZzdA
pjhcLqcgfpW5+5vaBHexf7iWgmJpMqTgFCkIkEDlUEPtdFdczmIcKXxk2nog6G2L
o36bdExhzsCAmSD58Zj5DIMQq+Pay8R2JmzWhMT0rw6y5JDMd7NeSGNXlXnlY51w
EhLT1liDwiDCTFwjunJkCOHvmSMB4PCwOebyw+BNII6RDTzAVqmKFFzznaiulSSR
CX0VV8Ti0HzxD5MOVF629DpsrYcOpY/37mo9LbQUVMfxjzIuG9zRyH1AvkKMS1yz
MkEUCnqirau1N3K4ZQBof2e8IMRvnxZsRuMmEHqPsFZoThWRqn5k0YTflcqupm72
8vALjwpJ0UPFszFg0O2UUraPcdlD91jiMkEhKOG1tvYxpBTCfz63qj17uJGC6hp0
VVTMMIHKaP8huxfF/N3RGWd7xz5QT2vQKa9phg9gNygeFoh5amTVzYuriK3v3CCI
8Q5ueZNq/lJDev704AKTpepahaYhvc7zXsk9u1UhyMTIhp/YB7I1TeetKGC1Bupm
kfUiMMsHuSvjXU8BkNobyTkLekEtuf1V4cO/s6ldOGSuehsiINmQJNTTn/MvKLj4
0N1vKVdUbuglYgx57VZ8MAjC7GhfXLqTpa9Rr8dKdctYslvdC4N9zu1p1A5U6Wji
wx7hlPQRKDmKEy4l+mU29AeyFqW0jfIdO3ljzeWlGpv31lO+L2l4MMWOnVsuCXYe
Yygaka8O9KyF+pQ0Pfy7bHgQ83XmNCt/Rda13H6fgBFNlOWF0vziPxKB0wYMoMqx
IPvVpAMGArdcPBLCN4X7vkEN7OzMFAPf5sCcKSDdtx49knHUTd+AIyS8RE69x6VW
2HI+QHX6OlyUUfavPXzktwLUVUowaRK73jG0xVxJrH0vW+rXXjNjmmSS8H8BEEie
tGptsRvVJnZOWkv6uEp24kgNBJwJ5fg4HsFkz36yjMi9szko9ZvTulmx/JqngASe
j6bUAbL61i9pwr5IIxeY/kNndWYde05uwYeSVC0++OtSA6V2HIAcGD9/k1s3lNwJ
K264dkNs+U+Mchtt06wqCs+bSJsCZHO81ItLBI02Xz5GCH1Y38Tn61z4d0UHYjWc
LG1ofoZZEurkrYVRQ4CVaGrcP/ob72dj27Bs/994cA42hTODq9V+Y3QKjdsSlscJ
DeRv6PnT3EsHlf9gm/iqqNnwuiarJMVJtHssHa257pv9c4jXDINxPjwPdVUY02+m
I7gsdX2bhCJCG9Flgums6yEgYB5HusWM+KV4vbHW9+u8BwQvDw9eztxbNcEpMfYe
yOTnpiGrPT+zr9tlklb8ha6LE+AZ9w6wKI+helQBQmWP3L+tf7EhFLuzRB8897YI
HtFXMbTdHaR9Fd+yGr/ZJN0nT+viGUD+rL/4g4aZPcCF4Vt25ludpimtYEcp2+7O
prRl9VRwK0a27R3xwLd09BEGtjUM8vZHmUmBPa8HQQos1JMPZRnhQbsaChO9UBGw
Gl6VOPP8Z7g81NDcoE95MaJgxhwwGTXcYur6HSnYmg1eNNDorzz6qeRX+Dfr3OBO
EQLbGTCkt2XH7IRIYzl4nqMpwHj/Th7aDy+8Vv+93h/efqk93Nb9fRCj4aw71Oco
05mX/Ja92mrPeWGEGJg2guSFOQjWPoEt0n1Eyhsjr3ljmIic5cBbtdseUFYTsu+6
/fsA3zZZ8fgCpAhA0yqK746cUciF56/Tlhd0MZ0AE3akvCfXTDc2h637koYDWY2r
CKiS5TqZahxjka+0v7p58DcMM4bs458KORXcPp+bGFwomzKVhb4SARMjHBiVL0V/
2XqETLB1raoYfJyvL9aCC/i7lNZkTrk6bSzP+X0cD5/3ESCsHBAk+wLaLYw6OKpz
Mbv/oHI0uXqGWjRE5c/DRkH6uHHYwXC5qHJqynwTMHbm99WhYUoewATxdu/TF8yp
eB+tbHLPYlQ5KAkNUhSLTXq3f62wXDiPSNLEAnIuQkxfwJZH3hCQoHS4meKozkcm
cur1H6hW09hpPeCZT2B+C0mKvwPUmT341IYoE97YRE6ft77QqVZErX8JmNKZz+LW
hhXwr1KItQB7sltThwzunn6OElfZrBDkrOJnx903Gr+qotwvruwHb4l14Fj4+OKC
cTWDV/4WcN0w6YZi6OTItEERtAxPmhRmm5jj1I6egj+OzkBTib3oBx5dKgGaycNf
1vX3uCNShp+KcjMfGgDPI7Nb/jJnI+Ea9iStTcwddc5bG313ovGlHA6XTDmBhITM
2JO+1fAazXaKwEjWiiHeDMvh2mLfJz/pW1DE4QwcTiL/e5pKblq1PSenyEef5Xaz
Wh4gJXxMp78bT6wZmCkyP89xild/f63cJ466zTQ9PUXBXh/ffJyyyicnL8fm2KCC
d36aoH5Xn7vhRxXDY87CMxgxW/Jol+MGTEjdUlB3agQv62A9G5bsiqaS2BTLwEgl
tc6VNlyYBhnpJjEKQaqcH0bF9NsTEcCaaw0+B5VUdWbSwQsTkxfx7xU9jSUM39BU
l9b7N7cyhox6M3bUXMU/DVXpTkAmiIMjKdNVyR7RjJQ25F4oaJhB8DrqA/1YwjNX
ZxyhdvePF/jXWl8dwM3eGYxBNcmuY1BYjeooWSmpUsvhdpJUrhiiiaZVNy22QFrE
XAONCKmQK/0pYL6nJhdnNkiRMmDcSLr9lNlvtF5u2mUTrvRvHfm8x58M1n0f9+55
C+IEFcIq9svslN2PAh0G4AwCRNtEKbfKwnIM3+64ZI/HvY/MeFjAk0APZQNn97JV
Idmg4MbNVcQKzF02GdQ1TYMP47DGyZhF3M4kFrSgREQXEHAhcbP0nR4AWfzg5Yln
oxvj5FYvfpLOLq1b07fj6UIyo1Q0WhnxJFUsm7TzwA7jz1dmiurOMj9N5ESweWpC
hdJY82GU3iS6mBZS+fApLzhYPWZwGNpehOnimfdGtghKZxd+9depLkoQrztou8fn
JvmluLxpj6lm9RfVrAR4mx/hu8q+P/fCmddCwBLLXxbrIpVp0hYMqoKKmqphlOPD
RVzk3LKEJ+zmc3P36/pPo0rnHI3v9ZYFhpBq6zOrdUzlfDUAVo5Jd5GtemWVLKtp
2+8lvnNTSt5LDh8F/K+bZZxjWpTxDNKey6ci+p2miV/gGk4W9uEod9WpvbSLgPoV
5i32e3qUzWGO7zy1VSS73mfCyQXDU5kUlo+hJYv+v5ehgvrMmmCPur+/kOO9OJNu
jNdtcq7XwZavQKAJir6y2MJ4iXL9eOlcbLryN68jxg6wJWWos7W7CH9P1JvlvaJ/
xiZgpgs/dPID62uf202olnPHKOS+iw1VqdrmdAgAfbvP5qrWB+T/r6tPI1cXDzkL
HIACNlMFnvGd22AJfui00VAQS02ubVK+Tai4nBzWWUNjPfbcFqFHsepbtEsExfe8
JL7YTeeo/2Av3jcKqLUMzQ4z0oJG2daYQdpkUmkcW8KcKB07FxxTtJyi4Lk2lQ/G
XgUbb+wkZkqVUy6+SkIyXqJicwTedvE6jjYfXZzrs+JbCKZWtapjsAZf7cTANeoK
JKXDZpHUOMdeAZg6g2jGcjC9kV8ZtqVIW0zLxFCrqXJDHMMux6H2watFJsOT26Ir
03Nn6LeOcBQAMPs1LKLLQj8eF/XpD/HoqgqBc8pYslU+S5NbXRt7HYTPnarZuE+l
OLdRfrQAN3sW+sIZyIfbfDVWESKbe0+vj1HutvWjM/vhern4ehsUCrxDz9b83bb1
t5DOpobc31/+sM/VSP9WOR3bXBk9HHGv8jeHeQVO16B8u5nSy0i2zLBDZVIQhJcS
ochRRL1q6xWBtgvRMXESSUv2nTNencG5BO/ALSvSjBGhUssQuNAHcFKes71InIgy
NgCWzu2nKqOke+BBOe8Z+e8M6OCT2TuYJwumeYzCp8bl7VT1caWiqnuSwu2heoVP
Q55DwVZaB3rPXFKenvL9iKa6/hiU4fJ41tsSojpj3Q4qJvPZMKEmQ4D/azzsuX2B
ow8Tw1GIBcpXTId5/WHNEPdx9wiFyg32VmZ9q85jK738YyyDi14RuR0jBCnQADyp
rzuZ0kWH2a5yDsePrMiNlh7FruCNxCEGWRfJEzGIOV+1qcW/OHRTIREWMtyCR+jT
9frq530nhU+YH99Sd6ZDJey+eZF8qLNFhjPg7memV7LpHLF1OlNXFaRna3ISKgyK
WMLQQAtQYO2UMXh8whEcBRIwdYwt6rtI+3rLas+Jx02VdWEtdew8U3QJmZhTUx2T
8hVQif1jmnh/V+ISgDc08kl82vCZcZhoXT7sujr/U821iZVweRAoYYFjaQAHevua
qoj0PsS+1INYjRRZlFxQ+ghWPT5x4vobFqJmwRDZ7dXPo9vG6vy0IdVMdQ6g3BHE
h//XRa2VXYWNjPA8tXxB8EzjF2B6WOO2DNQWms5bT43+dEKpynBdfWxOxftOnt3k
3doVE+EfksPtez05xF4opWxgotJHOpasxjXtJCsX4CaF/y5eAZFQBTyqu7lmSbXD
DgW/CJkYEznPqttQCbvzJ0GWYO8r1wIQUaYcY79KwuqeAcLkB10mMNrAdCeUXU4K
XNs10t0Zakns+rZxtTjzyzR39pMpV2EQGrrS/ak9W4AZwfHlY7he17jpkVcb6D/8
sZBRzUuGRimywe+TkkLksDkxm4+B/wKPnUzJA/+l2gddJ5Y+bAnkpnYIDbYH3hk2
vrXXsOF+r//yzM6TQ5vTSo2NmlD3cQABZ1lTy84tNmpQ5ihatOJ1I5W4BqaB6yZz
Wl94VY2gNWufnJ7b/xI6d0bwIf9Qls7jBGHnKMwGbkKErUgsFewo2ATKg0vF8UlJ
O6o0jX7mn9+MIDMz8aBbPlW9HWb+C4nEH4+6WM0ByPX6ukYUlUerpXRRTUkkWLHk
CB96rLWV5gEwqTtdVCrn3+mshYjLg/XmasoSgDxUOSdVOImevBf/SKVVDLqbwB6t
rOuezOAvRFbZ+golkiYLdo+STRGYV/gD+SN68wpvh92WpEd2F/peIpikfXpQvs6G
g5B8d+zi9NLk4C+t6AMcgfo3Jn2Gl0QJaSOTClljweUlYbyvb6Acrq7pnDz7sCyh
3uPfEnV8VktYbuQ3yw6xEl2Oexv93+VnxdjEE8dpjwPUhPi7bUQCmx5UZKlqsYWy
Bg6HYEc0huoetNgsTqzRAtJA3E5CyNBUgALgNyWf1uisAB0uYzYyv043zQERoACB
VgqNjpja5was/1PEw3hUwv2HX6jU2rncQ9hUb2keGSzVSad7PLsQx8rb52KOb7fp
W4AN3LrBtY4Ht+Qm8iqTEH8L0ZFmpKU6/rgqp5fkGKdokX24LblNVOxtEysgEXib
HzxMVHe6Li+d3qgq81QwPpGRjAZjknD0Ig0Dv/paIVKEtLAZBAsCa58PMRJxhHFi
RBvn8Ax/ZdW8WT/clry2S5IIcal3D/utiSca1YLqbtG2xTd6dbOcQjIJWZjVgTy7
1EbyxOASGyHJIY9T7QkW1HhmOf1Vnrr3xs/vTk10+uhEoXoZHgxdDrK8zaQKgt6T
ZCH9GL+/6hOpN5QQ+sF2OHDFS7ausop1c7cLkXlw4RFvoQxmf5y4iFLGVkrJkghz
QkIKTQySqSLBAa5P2tshX0CxUa2WnN9fdyv3GayMGKdda1JTbfXyGiucqChCG8DK
CiH/gpMUfcBSKuOAmJY4PBRGIbI6tYRT5N5X3uYklm3MYJ09A9f/FlYIXzV85ni0
kNFqOlb9S7leGsWvjmDeVu775MuA8Ys1EpZHz8nWzwgjdycEHbgwf1toIPuB95SK
rHpkQ8doarw/2HqRfVEi/zYoUgq3QYZiNvOQHT8lOWL5SBbebFrAfjqMYOJGn9Hf
iIGTtvly92gHNQDJQfC3+HcpnW0XKANydersUijeCnFQqExfNTCgJMs1uQkBZxiK
SDJe+Pi3r+1uXg9DxiA+eCB+9xL2bh6ZMA4W+Kh1DRRDjPF9g4DtOs8SOd+fAx0R
n6gUmXgGiJAHsaI7tU2HneW2ARNlJMrmXDMEnlY+AOHMLH+Pl7mm0j+kAJwza1/D
uHYgGdkAmk03zr+Hdv9UscWwa5ODJgR3mLAKXfoYg+3OtMHN+kiLW1uqXcj0o+IP
ks6CBfBb7smhfI5s/MgEkeA1x0CLd8VCKV2e5wi0e23/+2XpLaMbc69LRDTa/LG+
J3PqhoAaiyz4ntmBzFRtXFdIsZTHkEz3QB8pSkzwHDkQlb1JKBWlHxb78PgfWI1q
dzLaXbn/NebO+20x6UaJGmPI++wguQQVQi9Rjj/Pbf+hQbHaNdf4KkwiPq6z2egb
dFwlYc5hCe7gmkv9OZKZeJN0dRdKZXgS1ZcXsWCmZVCv1rzY6OUDRPqaaOUT1l20
s6Xy6saWNF5lGUi8dnjklUreUD2SPhR73XiiWPMzhyU9D/qstvs3rywdxW1w5U93
+nUxQweGk3/uya/gHmWT7jgG0wvWJYjM95qgwcqAcYlD7aOI9ErfM4wgsiPRQn7b
3dDesUaKhqiHw3oAhH/Vi+DCMjWG3fAF2iT16D7nfX/hZPTnCytwld+xBx4dmZsC
eCkQyskhgJUlTyxra+aRixPH51u1ICJsDbak4f+Q540MqaP9UOwUuGWNvvwmxPOT
N4XGEg62On1bVd8kF+a75SNojphQbapx8V9S+KPW3mvIq5GXRxZYQlgg8R7ISYub
3Eker8tLs2S0bsRhC9IIzrV3RgGyGX+//mz6m5MmHP1up702X6A7nGx1vQQMDD5C
1NEFFJJ0Ie0vPBopYA1vqsTUUo7R5GPIMiXx0okudfMgLHnIQ95MmVRFnwYLf33I
sEVtC5WQdoq4DmiZqejVcT+CJPgCsTXx64Zp9VyFiFr0OKVEzvuEAG7o8VbuEq49
DjmMy47o5PSVNa8rOlx60TuZZmwgT/mujQjiFAcV/gzn5N9PrE13WRhYb8UGUGCs
Hs1nmrala6J3zIW+pgaDC+LY3hk4VUCh5u78aZIup7N3AMb5+r9YcUHjorHpS/Yk
SgLTiO9VP5L2Jmi7maVSwdAiG18bIf22YkRZI1ILkczXV+1PRzCAka4N8CxBsppJ
mHaJ3Aaeif+2k8JuCpqKxR82kpNSpAO8LbdFxoQJU+tdywdFd0+Sx/xTj3I0hABh
PrPHaZ4FL8i1kIAHd1ix1BU/dm44cVhIgw9c1CiRIi0FHX3ngbVUnoGGd6+WCSYQ
ytw6XDXm4Sorxb36iMU1g607WYUjp9Cxzom/2e3JVok9cwocEHdqAqnkTf9Z4fGE
zZExbzQ7Y/t/g+vetCuzaIRVY7Xkhjm4i8U1iJzh+nrIDxRdUYV58ucnXm3yK9xJ
1Pvassl2RVajYnbm8F4fRB+O9IPd4TYjYCPm9Lgq6pcAo6yNwEtc5uvT+iU8KLRB
uLhHgAHq8NIL1gxDKQgupFwI34A3XRGEFOiakibIo7DIDWkXwCSXs5+dqRh6Vko+
3OBEUA+ynqQlWEEr5Uj76c7zaMksnXPjgrowLQ1HZVL4Hgx8MbaP/kXbQiqzplYs
itWHv3b6gg2xNoiksQPUntQUCoh9jfu0sfBnWmeA8kFg5wBb7X6ElvEb4TCT/GZS
DIsfENn7IFObnasZOZkosKUFWaLzCwicWammYniyMoaacHBZ+VKsb4bqrCHeg5dO
19bcEVldfmFM3mqhe6Xk0aMxJwl7CdlP5QiDtpntmQbgOe5HRl/ZCeHEHb3n5EHm
JEpOw7dZFuIZGxxx0/ao2T1XWbityBVKiAmuu1ephPrdNpKFihUsgraKOKrboJSP
Tp0efyNyzLHA/zkz9tURTO4uelKdsG4rrnYwTFyZPyr3OOWGMvbbPeMGeSC60Mvm
hI5lG9mvIqHeEua4SS0O9FQQ/DpivsekZkWwW3+KFZwOURfGjdFAaAEea1xkWyBj
5hn+j9QvZ7l8FRoH1dflD4RWeAPczLRKJGoMR2xJ6DYRdSuCdT/FE/flGsewMy8E
zvRZdXsZpDyIkR/lyO7kcM/YO2iYXITOrDNZzX2T3vy0CSVYNQ2YzMhnRztowOX7
USG3lxA4D04fIGG716EC30QLonWvKnBmLNkVc1+UqSHbQGxUmkelXjtq1py+81nt
GQtJV/Uy3u8fBFH1hcq+tACCeRrwzvem920v0peVf/Lmvs8cMuadiEpbdXMCr0fH
5R2z2S2G3nrNqWPS3E3ascMqsyuSHkz+x+2hX6aQp9B8lLsIblmQ+e35uPFt6liH
zFj2eG4DT53Xgvzw6cF16NGiPGp1vJ65bOvA2Ryq1WFGGkX3AK7cAeA6YWQpnWcz
RScLtdu6WjH9/nQQFZf0aBKXcXxmrN8RShMNM3JBroLIsaPWJylkES0lVfBQZD4d
gMlkrHKecsPIfhu+2419gQzudo01Q4LY6EPDlSqH8jH7zH4myuxcpPI5DSN1gd4p
vbAaQ+zz2zuXhik6j13K2L6YHo797X2wgVctqIzcfQtaBm1ysVmE0fYSd6YiTfLQ
FlNWQB7IOaydYOUm53USkUEGOMzN0bECEEV/+Kjq6qitLtgv35UgjNbKUYHydey9
PTn8fmhdIw8j9d/DZ/6wrqLhpZGLAstemeVUqPRrL01qCzAmy+oG62c+JAMUiE60
zPOEgolsx0PQMe7uPbHrKSczt8LHHbOVsPn//bwEKZ6YNHYgs8VPP44hxYUpgbZm
bqesn+A9iQG+YZmavsOiebn/c7N7X+Zc8cIPsR3GnW46QgYkP9LZEZ7DqbSgewWO
Gp0enQB+10k9d9dXvKbm++1hN5OMDhvo9/Qn71qshqjN7/qYBixtP9a0tGvL5Wui
NYI4ILvu+73AmfFVWjL2e8aV2JaIbPGvHJ2THxb5NwDpnmGONeaRfwQcmqCsKR4r
fJiPXJn3WUnIKYhZTBzlja9erIAJL9Ab9rTByyTqLaGIq/7i0ibv3jBzHksn7Bdc
2tJwDQSOA984udEhC85BWo/8CV1Sbmgkh24v+XIWZHuw1o6+8K2vUF+d7hrCmLNM
2zgVxN+DVoobcamtxN5DzkJAvMZngxFgJKVVRr5DrMrAHEmmUhST4hbol8g8C6g5
8xaiREm5b/HZDXNqPD8KT+zidjZMPHLBRUWO9X7JiH8eBDbLkMnic9n/phWZoTUk
65irOVh+XOrYwUxhqND++npnn4wbROmZaNyQzS8rbX9gYlTBdf3E/7Chvl5ipRnz
kgk0/fAEZukYSQZ+mw+d+rl8wj6KJ3clga76RRLrZcirffkM96VY9dsDz1yRpaDs
v0eBjvzzk8MTJdWeT9JpKY8BJdBDdsAuQTJLovHqadNAQnX6YeWkfPTkEhEJ/sRa
eZ8mM/Iw+5L3kjE2TYsE5fMJdlBakV/H2DBv3RJUcJiayWvlYKhhQKHRSln1QQ7p
DMxQgyFx8i9ZqJ+44a0OpxzrcFp3DCaO+ttmMmHLh3DDOURvQkJQ3JpFBfulXZph
3kv8R1jm3UpLN/6aJEGNqBGYvlPyUkqegr0cpPIh4nTpBA2jrWzOtUJIP+BILZ63
LHCxzMOUa3r+3GdZUuQ7eHWr+eDACU5YbJfYYEL9QjxOTbqtnLeMba9BpT8ArBfM
8bnYWgJkEfuC/8PaGMgdd4rBEsb29wF1uE4JB/wlfYqszXZjWsAvfhy+NxqvDDcQ
nl+8h34XcoP58kj4WuQ94k8bXm1LbKRfSa/U+8XwXssoyTixW4idmsSN05UlzF40
+lWLWG/fdu3nfo1n9FU9cCe2Maz2kZ8SemizsFqaqjN5+vWMWhszKBPpOAll9jS0
fwuf3yaL9VVUOGlel2ssFX3piH6HLXSpDOiWppEorR6XpV/rBz550QYRPv6Ac+pF
rMITePnSr6nLp1i2zYIC4MyKH//1jtRuFzkdzLCbSVrX/oOTwSMG2mi4jy6lyS2V
hpUEopEtCmDlKH0Lgc8JFZTcChtWBA3GPl4ayQbTcl+T4ib+Rx0XWiGB16gbMv6X
A37C1DHTD6yfYE7hbumkGidUaO6ah9rxRsl3do4wa3JPrScbf0nOi/YEvNL0KJTV
6KGSCIsRR20WxroKs4GRBMh3mNFKjdAuz1tek9Jc50TUxcEGoljLJem+YBNKcmLb
Z9O6F5kmb/URbGTqjhl7s2Ol+Rw/SHdxMNl0bu94u+PsWCKsYZCwsmVcdVzOY9o9
rZp3k3c/y+dUaPjmUdwmKmzIFwZ38htnk3IldZDaI8yrXcmNjZuVtetnVCPQS3Ee
Gwm+rnjz3pFzl4uXjs9i2bfjM8Sq4wgTPM4pLhr8Ect+NHwBT/FwqZqXbNH3UPe9
kTDvF+bBocuIhbJXw398wU8JkT6SGul8i4z1c1kRqQ3NInMUyVYr3/Cm1yLygsjq
+nLuNOMkvfNd6GNPxDmYFVLCW+F0Sf2MwsfSeoFmvfg8t/a4JwUBAH/eHlmzNO0P
gV3tJx53pWqzRBPd3aYs9UE6WARCkprb2NnK6Q+L+ZuBLpCHo2RIP10hhwdr4tAU
PMOMP6ZM65hezJ0s8DbcYk6sxiOUulA3UF3L/uk8+fnSK47iJH+dPSjRW4IbokJN
+ahHEsLVpKo9QprGAcvC8sTuztbx10gw6U/XxYZNhQSGYvGk9nFEtvBB6Ray6xtx
burci0EFtprnhwJVQ+HvwwNLb2LfH81YQ3WeV7JxUDn5y5BhRQ1KyTWuUAQIua5w
PuY9gnRm9w4WEm8GEz5Ci/Eof8DCERM2TI/YqoTaOHPR9rKXpjWCa4nchRhLlToa
U6TVta/RB6jYa2iPaLGdaULssIrZMl8BtFFU91GUp3zXqju7dcN6nu5ihIuEJ/RZ
2wH0VVoalx+SqCP/68msL98taG9b3SmRvuUSOnW7d60QXU/yEUZ20OaVTUzXE4wX
4ak3E37YMFBEzX8/PSnPvM310N2OIoP56vNmirXnL/rQwF3HkYbGh3U0yQWWFsRZ
4nf1ShIz5PeXGIvNwCAnbO3m1E3SYxK4mZ2pFc2egrHV8QrrOh+4spgaOXgjWvFz
s/d3jMm2UUkuoC8xe3NjO/RUctWsw/kcNHK/BCFwhmmMtKVvHApdsZdfQReSTMRL
RS/wXcAH44bZU1kPg425Y4iJuvkLk5IKvpKWx7xh6Fxt5gxhqb09GKp/APMhqJdJ
P/Oit2M9xMJOTdXlEBdPkcpXOICHOpK9/VkX1jQMShFCaxKzx0zEE/a+5TtjsyKG
TsnScfVQpo+gD1LqNcvdEidywlgIBwHEgSfB09vxAfLsBu6xbLlibmb/eTtEzovR
ALjVoi8w1kjlIwaERh1OdlMjdHAmx7D1WwZm0p7F+TLHW4yUpbXy7VCQ7mIoiI41
jvuDsZrAZusBz4xPsiddAS2wzloMCK5Ed9BlrzwbbUpE7D1m0seLTQudvOO3pCV6
RQ28r5npgj25wZeb79J8f19BnR/A/rQVuRShkj5j0wrrG1UKCDFIQfymAU95zMEW
q6Qfa+XAjtGl1o+FZJnBXtXGMPh0LI8o3wsPPPc4f7m0D9yDBvMhQkjA3owFyi1K
rUQc3QjrOduTkdr24jDJU6ggb71/7rmLojqM50w/Slp4wtt3f3AlQsPfqpAcOsPj
UjvhFS/MGf1qC/oCgo+eT6ZHp2D81tlialDOPtD3JT1mCEEle4AGiWPemugFi7K2
blDMleiVZl4KvYQbDC1JYXE1GIw6rsLw/MoAxaaYYMQxW+snBB/wz167jvikt/6+
YcERC4H21+iThUjEpFBK/AQ+MKUaSbmsESRjrmI4y0qdto49ShCuulY3HYfxMel8
H5hBobLwzapwCheS2m0A5qPLwRmFGwt5HKv/UHvKRniv2doPY7s+GNtIintR6qyo
uQPW0ibzMnofzTnAiPdHSFFpwEO1wISZQQtlgsqA3cVqRXs4gHx4tXtgFg7kJq4O
27y4ZAQn1pn2TaRnSJ29MFr+XFVWUEGvr2k9dzw8l7u9/qvBHrI3u5YYclzNaQes
t5VQuXxp9ME1TQg6CDoDs1JicLb80i5fA8411UDfNTB2hHoYIp/SBici/Xix2frj
/v4u0+BDOA0yQ7KUSZWUgy9R/86m+ueCjx71In4ynADwXvitZJlmKiCVqM7czstZ
GcOa+zBYCSdNUrI6LSRkZ4HPIZKLeMJHsEeYWoDzkY1cx8t8g7Q/U4sFFnmbx1Jl
Uj/IuHxi+/dV9a4ZNACEWtL/CHRJVPI/nS1zwYqf4aVcIeX/hrkcbedGQB6wSIlh
R1fq/oQXxiD1fF2TXjfOU19/WByEenB3F+5olt+bVJK6Ocqm/5Okxq6omelhmeN/
ZmxKMumUmbubLCK78rW2+2yr8gghCgjbn86e0uzDg94+VuZ3oqYeVorUGCruFn9w
EN5bgGhGybw2T7h/nktmMaX3Lz7OYMIPbjvkO5qGMwkvuosx215Xqu5Jl3nDNaoa
bemx+pOz3PRJCf3/BObsHke82miiIFLiISYVz9N3ElLRKAMywiyYBhkXemaMyPMP
fwFpn0dba8eSnxCdHsGrDnVRIY/qG9JJUqfCeWvcDLPchvWtIVJ5ls72djIaexzI
45tTHb6wl4GfWI4WsYuOVcOoZYPRfpfRkpF+bXvxrQVLQ50uUeQ1t+JB73PEdBXo
qaIkzUU5ina1qDx+h34OVUnCOCI8X6UQ+DAVOXMv76sgepu9f/cjweucm8drgICe
/1FnPFGFT35LNWqzBdrLCMUd7ttw/6tVtulWNb6OGmRS3FRCDB20aFre0TY6aosO
M5dNhA+iYGJk1HWH2AtMqQHGWqsx8LId9ennLwkxMrFcX1ADGdJrsIpd63SlTlvZ
T6bLkhYQrecJzzOvJtyXPQXjGCseocCPzFVOvTZl7qGkEyef4LK3uSazOaKz+JEA
RxEPM+cwbSzAt/SNtGl88QmPVhZTCapf0iEXqXM9zEe0EokoTdGbF+gVzWxvTVlz
Xsot4aa241rxrTF+v92COYAIhup64zT2nLxmpyFm/y2452vC3pPydCX6J+z35yzK
+oxNOoryZ5YuzCmEzXUcYI18MrSGjyV2pDLDqlA0i9Kvkbu3i6uLsKPXAl7mok3V
QXmK25vt1CKphW+nFxFeqlKOR17xZZlHMRl8WM5+EdCDG/8aFm5jWt78C+pF+8vX
iBbn9SNeFuvFtytNf1ObusAuHD2f8D/n9m9rAiGxjU/KY5H6tLGGHCNNIu6YBeUa
I1r/SaVbvVSg8y+CATeddlQ8pQfVnsPajxGzwAJpXyKRM1+UIiyRLHSVCSYACXgc
Dw80/6qi+et+JJUtAFWi9RDRbjU9JT3m91XRBfoi1iiYopUb05qVe1deNQt/0TG4
u6PVGu2n26xaqeMqzwFAn/CgOHdQXfmFo3lBn+GDVvNY0ihyAaoYAKHN3s7g35IG
bh490RE8FEJM/NEw/2DNEYguu3k3C/dDrqv6wu+kze8OZC/SBk2pxy6WJ+8FcBHC
ZbeeZ+Y1kEQ6SXug0dGwNUsCKJSkjU/HoiTWBSxKaPpMHdCeV3wegBeHo+EkyzTQ
fEcf2txKlqINA73Ctx7eRDnhEeC4YY84wZ0HfwI5XL44WmoGd5hKZLjs7shlEp7i
/EMPmSVZov8VMy8k7KlotYtDy6N3guvbJq/AN1UEcLYEl5gLgMFbZdnGQqltFEVq
r/l84FcVUjlOqLJhMgkzgDDlp1+wrq9eZf3NV4nFYLhSVVm+P7ps/aOAnU4h05RM
g1RBNKZ0EDtN0EXZ1AWD1zKbRBvAyxkZHb1LowkIpqAdhKT7MtsmwG4C5nEIthSi
6wrAQCYlRVVIbOsZtJfxcs8nXveSQIooNMc2LN+5pqUfyoelXrCHMGMGZ+vSQmT0
HYB2/jE0PDVgOW1GZDVJWL5pIAD6boS/j53PygN62kazUGGH+GHufNDSZ3oU6RGV
8X/99ejiS2BAqeA6M2kKJxwyAg1KfoNSInBk4hzXfXJqKGs+QYKd2PZ+7mXesGf0
mWjDd04Q9qlktBmI5uMjD6htxj17GgpkPOzMxs/biTQj5aFO9Unr0+9I8qlcTbb0
o2DJW88VULo6aCGDjVpGMiLY2wPaD+Azk8CZe+7KxgS/KkKrUXljHa+CJNzuHysm
HBy/KTr9JQsCSJ4PD4w6I6mLhd2u8IGr8AaXmfpw/7Ytb7aDd1RtkrtyxQobE7MT
dHQG2I34hjUPdD3iJFMtN4M146Uf0927MdayDJx5OARjnOP8Q46ICR87EQeP64QW
Q8mQfYS76edziAd3r8En1OIWUK6BZNEwL3nxXu9wOHi+hpkF5DJmHYf7c+E3BU0K
0StoOHPllxk9S4f9a8mHZWEDbkohhP3qbiruw5QyXJj74vkbBkTu6udrmoA2yh7t
9S+UX3H6mODB5XqHx0iuzyZrJUC06wDhgIzN9+2Ce8aCRW0sBg5m8dnvsZdOf+L6
PGz/9j7CTLZn4/I9dS9s4Fbxi9pFpZhaxkEo5BSQJ3wfZlFvfAVE9mBgi/9zWFq2
UShXlWcYD4vApQNYqoWl9Fi7OowntubA29abnyuPHdyKF7IUSQkpv71D8q8ErAII
o+KmVjsrTnFk6gX6cRGpD7ati8FJ/WpB4AtN3UnNoZsfXB/DtKuXC0EISQTP6sdB
chz9jglkqu3Nce7oZxdca0ngProrWWtvsDP52AIpClOtIO8G6XiANA+Rxy0ZLFvv
8UKFcJuYkvhxngMo4bOOCaEtLQXS/Kli7tYQU4988Ry8K9/LwJMhIjc/JlD2S21u
9h5JW1npNaQR9BflXxsS8pIpm/bQcM9oNKd5hvV4GlZgx3i8BNvE0mg/UYFhVkMu
ltMcIIek0wxEs2UquMa6jZwKhnHO11N6PjJYQfRbwoOxF2fmiwU4W0DK1/jxyDjD
PhV9A5YkaCHl+jLRKhuVIqRa18PCbCObCUcRtt/TyYvWVdY3IMS3ExJnmc9U9dPS
Z63P77xOVT+hwSWB65G3CBkeYi+c928oEcvC8YjvCrmq3+JW124IJYFCjSoC1/Ov
uEcZsviI8ZNOIYme8GdUCrgpotoBG9fOQl19kVv3GEOcFtzoCfiq14fe/Ri/uG+9
ARQFRO1qRbqUF4WJxX2q1sp93rG2aWGTMpIdpcBP/kJDED1UsRVzmWPEeby/5zdr
4sHiHtPiycTyifqaEXMSU8UWuWKcoBwonRguwK5/dnWR7MC9lynMiKTPFrMroDWf
1+SSCtyEQjLHBhCuZoPyeE9Ifta0bH5HAfawGTJLcZm9K9AbkdqWjj20UbSD6ida
NCPyBhcoxAhgxKCj/Bz50KaWAHhrFBD6QssUguaWah8j5k9Ribeo4bUPbyKRZSvJ
SCf+g9kdR5M8vpsxTs1zUs9SfQwzNJc7NmOvB1WGH7T8c1Prg0vca8zpsP4mP2Sh
RuKQ7aNPGNpQHYwiaCw2zqXfNec+mwQ46yyK4qxxd2tET2+awbUJlfVMOmSgHl/+
QoEK/1YMgUWsbtRULV6e2zzSMmD+KdH3nA9NlT/aJFU62Ymwfs6StBZIdfM3JdhZ
8visoi0PT0lQ+M6HaUpRokkbP98dpTGN63QY0OTdeUR135ga/YDbGdf/TMkhdxXJ
saZsy9MwsnptLjTwKeR2gncsaC7rbfTemR1HXL+ae7I5qLofgF55Ty88QUAwk3jg
Iseb2Oa/Mvl5Su5OMdk2IdFoC1GzCoquq7ewGgxeeuZvVTC/qptfkonVlIDJSls5
hACbsNyCdXo4+Z0aENtPc6lhuhRwaNuCJFck/wUo0QTHiWnxJoLKbfND1EdB0hJg
1BqCMFQJG2b77pxOsOS/EfYAyL4UKp7F3LxR4yeSEym9xNgSVhogm4eHShqoZXq+
hBIR/vNuBUIkBgM0XzbrntT2+7eIVtxUxr3BFH3xL6QEECgq1ahLX9uh1vs3CVJ+
HvZBsxIM42TJwQ+FHTQf/F1VY2gHAhsaTDQvCuFQrM9AUC7EjZtz/2kY1iDCnTof
SJtOcM1ixEEp88rR9RfvzcRJ8mjRF7puW+gcaZZe56WrC9PSitkFTfdSXbvb+kpT
4Klv5Oys3cFw9M/fRXc5CWBzt19MhoXaNKTheoQESvGFCFesy/oNJraR5g++0EHF
uv1SQZ04i2hYiJpSqiNo4ApS9bzKzG5wTHn2LGUJhPkOBQkbnnd+JOIl/H0BvQf4
Fck6dnDzUvuaZQWVc5K1H7ym7V/TpjwSOalx6KgzLl6eE7qAhqnV5FxCzgUrjSUu
ylvPTXjqQb6d8846UiCts1v4U6SdOPKr0F9UquUM6y/vSCKNhZeUs1eemWuGNzZx
VZFHUyyf26NSexlTSnoYQk4cRJqEHjeX1ohXQ0Ny5s/bZ3nIZvjCSjMCTd5mWj17
oBHVo6oP/tR7IrkMcf7HYO4AheJe4iJaVsNNcP99WSNGihEK4N/yXNJ48QKcWK2l
Q28rE86YtQoqJ5tvSVW7shPUpfCIMGUrwsoiZnQBFcfRxPH9zybu/hbPRQ+sgSg9
Ya3m9Z+b7oJ+UBWJlnHdxxus+QBVceewy6bZLbqDLh73cMaRYw69GjnUlooJV7bj
H8giB2w2aINvEoBqP0v0eJCNQe7M5c79ueuduFgEefsTefVnpWxrO5wbbBwS/Ekc
Ss6lC5sUtRj6tHpc2S8StX52eYeHsi+5QwsOwA8dx9C/JGTuAozpKCgW1VOwKy6x
63EMxo4/wjUGr1WkZhX7a/3txxg2hht9TUcm8EGADUP6t8SUCZTfiIleyXRtPipw
eQRiUkMbjzVr6xUZlriyKB2QS2XQgAayVcmXAgwNuxvdPComLqNpUN84LaNaW35O
Tkn2dbrhU53wObX6jFndg0IVm2wxnJjYilzC+pLxgX3pla0jwY/VmHa0TODd57vG
UfyEqrJ1ALJeT0Fdi6ldS/UyxAWWmJ8RiTFgxmxvMt3ezyeFc1n3AvQQVZLeJieI
lKZmuxHEEGhPGs40IF12mNtCuYQrQgC94QtCw81XGtv/ajGXnDdfKc39hBzR0ySl
9GXP18ZACyMRJoptBWaZa0HWEgMFsZvBfnqWFdHiE/EDhdJLGYnAAwXOU34vcqGL
ZepH+Hw16GiG2fd5LHxt2XnGIGumZ+E8Bf1ZRHdM6v7T3Ywg3uiAhs9EgU7SJFRJ
XnlkPRUoL8R9y/fw987GTvbzC/FjgxFJiKr3Zx7ivTbBXDw4pCAmr/LCqjB3OuBj
PnqsRqEPcvCJX0tMMyxLFdpjXcq4bJuIbYCUsIGxHt8hcz72X+eHYcvAh1I7xAp0
uAwOxFJr9H+6JM7FQO+mgHua6+ODp98x8RC5BbkfK1/LM5Ox2atJQiPZwPK4mZPX
Lse8kFMpEuWPISWO1cIn2djyGJdZtWOSrNhMsAkCxNq6c29TKC8nub27CqiLYzGT
TDLkW/TinVuRqijpJ4Xh16+bxu7YLLP1NMgNlbgaHbQWAZiNMzJfgzsGfsPvDk/C
30FPKYd2IZwDOSqkSA+slf3hy3jqSfnAiC+ZfUstRrKkS3PJoaeuzUoAOL3Scal4
SDpO3xLWUZySvfqdJKmwFUg3aY2lDVkgS9HJF2YDtRNdvg8B9XkhdXQqXSwS5Ofn
9d1AHSdeQYVRdWGf3FTNbN24onGflRhc2x4/MOMcmrw7zCuFCkeFArIex1DxvOAs
qeozXjGteALksciGzj9Pk/aPtHzizYmzT+1VfqcZtTj77XC1SbrPpsHUN0u/R5BT
nh3G4J4kcKI9O751GxFDotVhLs+j1TfIe1iWRx3OlgdIdQFszT2SE9Po/8guKlkO
Amwr/Mh9sFnMzBX+GDPhEzwSbIwD4DWpNayBa724nPGfH+27puPmwdieVJ/r+b2q
yqcy2OZVAr2FsC5A5qbmodoaDPTBmfbsKSOv40oTqBNH8GCzkOrZ2oJ3eDWX2Sdc
UCs4xuEJrn/dk3RVoTRyMy5IvVs/c4K/41iawnbFNoIZmheRB7qFrBrI5GKcymvA
+sSXLxkqPXx/TA4YIwri59dJQSVqmy0XANpFRUFbHeUI9g3Lub2kgJIxWkp+x5oi
ozT0xUzt4dSrGadlAsnnNDhQ/Szshefak6Fo+RDkIt4N0u4NSXdQn7GzjW+4lEi3
OdyrAfN1ef9RbiXhYxPGpjWw4Ngyl9BGOlXX1a/VXC2edz6062onJPQ0HiX/NuG/
BegD3zDnp5hvuHUMpASMEEevMEALibcUZTAQ6on9BLMb/pJxpjgcVYNxIiZfHkNx
cEocyCd20KdIKBuk8kO6sefYIBElHq+qTKIxxxcT3n9d4hmwhfh0LotYxNalhYd7
k0J+g14y2via7YaSaMc58v1Y7A2HscowsICjxCcw0jN7Qkvq4p++QOjjI2b6yfpW
KxpfDL/s18RxhBDHzOVHIc+/t/qKJOfZFqiu0TzZmM5Pe1FrE7OfO/YOa71wiqyk
uYUZqDjbHTx+PtJ/BPQU33JduHtGQDCmxh3fDAh4Qt+DDsebHQ0yFQn0a57InqdR
fIzhRX8hFxC+DZX4AEB9SxsqakgPeruVgQFusBAaCcddifcFPlCAyokpA5xVYH5W
hlEVsKxuLQpihHDOgA0tbx574SNhnDdoeI0v/cZcs5gE2nwE56inGOQ/YCNM00HO
NDp28MjtF1w3GMtZb//hbF1tneTMGbOIus7q3reE4oRLi02TLi1Ba4vTl9CtGWUR
RziFp33xhMCddo3AZeEo1f7L3/khYxlBBpWv6l5ZHDyL82j1Nvcl2sGq7aXb9D1s
T3kFOn4ucPbkqLI/HSHypllr2QrzX+bDkSwkY2WYPhU90joUt0j0UZ5IOLpwncHs
J6/R3zkRI09Xr/e8nhaRYiesppjTk8vRInHSE0WL1Ayc2rILXynbupuQG9IvQItr
L5Q7z0Juu8Ymv7iQkaFgsf1PGXRCm55czJJHstW2wFgv0u6BQtWB3ddyntb1RKbl
YiKIeOipemc+UpAq0Gj1E5BOybKGwd13qJ9W0nm0ZfdFPORxq2N4MVQa+u1RjYhx
YnwjqH35ivNFADyqwg9sGrp4AsU6t/3hKcy3lHJr83LeUb59PSVZIBLaz400BZaO
XqV4vSmUhzXd4+m/wVasea2Y+wsp2Ww4ZiXEM6/xFkmFmNL2ySVCAY2lK+IbFSHK
eGgolPiKZoRySiUyBPEh6mCAN6tvZ9mdq9146sRbigeQcmcbEvRK68uyRLqRXYMX
IVhqaSRRSO0jQMNAtp0uBqnnEJyUAN0q48GSbeysW7yMd+WQ4s2g+C2HJ6hpW7Jj
a0An9LOrvjdwuK+kp+k85/wJHvbXCYqUa6LylyRGaMC+ikGBXHSIJ44odpxEXnsI
raCpsR47/2kT0YltICdLBjqMxiPuhMkcPrZCJir75JLrt8mH1vRghrtFBhf8bDIp
DjbnU7HrgAiIRdG/LjniHmlvJMuf6JbD7/S1VcAAP+Sh4zLCwcWAv25+y9plUZCA
Mj9e79utM1HFtB5bUTimZFOJ1Pbipjs+wnVqyLSQv472aeETDbwCewVb/mmi39nF
0Z/JxH5hRKC5Pg+g8t8+7Hd4Ec+KnmFs/MSKK4tqeNR28sBC7xNIhVigMbGWorf9
BNe1MmsMX7Wl1M2AHSj63z7TwiqJG83ULjN17A1zikbv6gV+op6g9dEDPODb9Cdw
8h4eB7wKBYnRfqyaZf6k0VzYNbG1l5G1aDgCOHjF3ih5gMPN1s/FoNQQ7dAIG0Pu
/2kh2oEOsa//p//VBrIDSfiu2M1KuXR/JNeENEHUhNygftrfbgDXfU69Xk9NAoQC
BztrD68BzEZuvbFVV5d7gQly3XiII7hRlpOQ87jZRJh+6Fl/KM/aNrg3o093uLYs
JYNuLZ6dwW2rfDiOhR1RfaZvBxIyD3L0O4b5SUijoc6FB7pF4Nf4T00Gukk2Y0SQ
vVMPjr28yau7icnE9mwaAAx2iNSG/qaEhgvHaAdNRMgxI4+98kr6IhhOXz7KI7kN
a030BvBvfbsj3wvwmNh8unH3lLJS42EmCN+OsBMCqwyfKfU22TLTB9gCGDD7OZ4r
lSjNVpoKqRtPambMDZPoYZboY2BKKVuud87jyC+u/cN6JMcMwK+9R/Z6yO/28H0F
lmPXnyegBGzNHxNAZVuMd7h0kboaKdRwOWqP4k3zH/bhpatAy1eN2xnl9ml7frqe
c0CCJXLeJcqvxuNzUdEudHrkqDzOPyRbovmCDMv26SnLDfeiy0aKpfAYvP1ed7vZ
FoUZOtQRA7nq1PH6U4qp53hCUGxt1nrlnUL7DBYD9f6Iy1Ne+qh3n3chc7kirnvh
HRNM7aHVgtWhDIAFdtvdWrx+J5HN1pi0+lKVakMIfhI1JJYqEm0EsLlf0fza+zIi
M1CRmWeqI03cqbeoU16FvObHx1gQNYnHotGZFAmI0d7uR1KJ17wBTMlswm/LjT0S
jw1FU3shq5LB1WqmeBxUpcCTc4tNveUmZpojR67BST396BiaIXtfNepAuzwpn19x
fd7ItzjnCs6i/v8FlVzgIeTu4gPx9gcMnim4FPxjoGOly/alKPgPYANOpk3SIPYh
FKbIYi0JbHQw/aiDNYAwje5w2rZ2FxZ60R37kcjAC+mCUhNQ2teBsEsnBbbRA8Po
bpARPrvPeHdMLNOS1WEuUvjMaQtjRyECZ66JCaUV/RC/fmPTDgaIcoFOQe7TMia2
GlaLMmcynDYW4x6p1lgyjOdoEghmnePCZA9KK1IGCBvO0ariPoKjFNJebpm+vUdI
6cm96QvcqeC7A8fUtnIjHN0UpJvhEQF0YBjBlYkfMN+d11/PLRrttl+e0cm4oBxQ
J0PPuAF2d9lX7TP81zcYk74Wf2LE6BkSlkqmiZ8QOuNpqy0jEIPCXEhfj8UCImex
47WPMzxEIBZdPhTycgniUBwN/ezn3avy/E6Kat+KRFGR752c20oe5qC1ukZG6Xm4
SKosRMMyMWX21i+xjq7P5ljS2SVrRo3e8+TimF8i1WKpmMwBcyMnfr1S1P87j57Q
xTV4Lbj5jkcEgTRI/Np4cYNYgN1xICvOHp52GrI7yKf//ispiqqB1pPVIG3PsInb
FjtUmvZvTuK67sklQEb6NZR8xCVzcU1pCjVnNZ8x7BL+eJH5AXZpFcz5MbKF4dHn
VFjwnuZ5bXuutBPe5SGSJfhM1T/4WtrvOihlVHpjq+JiyGALWL9DIXqACXVBzEjW
TAlsv99LvB35R40RqA+Zd9XbGM7xC+qaUqVMQQvPZlbt16L3OcH0QYmdG/cgTVzC
gCRQBA+Z+pGqbE8UXu22b7Ki92KlOVbjXyvc09mqJyGsy40ZygVU13Cx/dMr62aQ
GAobxFVwXzmJmdPWeLoAUBHTN6W1IlRWlW8DpToinDVlI5WBSc1e7VzgU0OX4IW7
KxxSynJdZvflqNqtus24nARVeiwlLosK02/HVYMMdsHr40XBrZ60l7YIS8A9i1ks
LBLQRxFkLuFEKK3LWUv+oF1woUWKqpL+pYrW69dmcfczxyoGHhGjbw8v6rtyoEQ3
dO6aAKJFLrbnPAarrOxjJjp2nW5Nt/IEgWK03SrD/X0vetiJRG8nvQRlgV0CQP2Z
CWBmGKXTFalRRdWN5NsLKhlGZv9DQK6JGvcfrWtmSB74Cu8BEl1+LXPidiRmUDyM
t+8GBD3E4pJSUCOmwmJPhsdztzE/h23kPWNhkjAobREBPT2IhUNuuO7MYMfvDokc
zbqQP2nwwhUkIuF/xvQPskq8pkrJn2xHU/wG4b6MFRKUqKluNmLA/sQr4gb54c6f
0/xnb+aTQeTl2zSJYKj4ZOMWuQMCu8KCi8+aQHrH0JMWiCYhtguRRPDdphbW0jGc
ImcF4ukv5wzQalwN76s/Idfw20ypugbwLnpzlqsGqq63JoUC5LnyZqyf+FsEEnAZ
e8RqNosKnkV2GUYo3vRcUX2oE+iTlQx+mDmuuU+nByzhQNjJXihGBUyULC+te0mx
TyLp/Pt3TH2HWlowqNDoxOmNiP7psjfzqmZWl2PW9ZCTbQ2/LBovvZas0y30eOPd
oCj05ZKbDkU4A3TzvLfl5J++itn7IlBBhFvTFVqiqacoiTJ/K91OnzA2s5kFwn7R
YatHww6rlTrwYLNmiW2z1NBy8bQnmGOPzesY7FHisQIVT2ogCrLHh18XTPISt1x/
yPlCri9n0XcBDIGVbhAKMwYcB0H5Kof4KLztUNyaIXLCp/KobyKWhG8K2YSlWFiB
4nSVm3MVaq+uxa/2pG037mF9jAmirrGXSo6zb12iFgXGMQ+Ya6NTKrwPa1i919Ob
HSKi5uozJF8ON4nyeKZ8V2NTqUW3LouR3IoAu+hf2ASQFB4XOciQDTo2ByOgjVhP
JVhluXZkCes0dEJDS6y8EDGhhiM9irWQT5tSET03SV5ckhTylsKkcU+hX9cuVLXX
DBmr9XZwVKmOD2OV82yN+1nQy2O1j8d2v6hJ8dBf6NVJ1/zhLDcwjlH4MoKnGODM
hnAm2+26zrS+yKykwfbEimsFW2Qd2Ms/qw0kr3zhn1TpYSekSJuz0/AsX88ONPAB
WLVm3uWqMpCtApwp7t9psc3wFOKhyqb92jFgFVdPjcwn64uDQ+D0P8zV3RKvyBKm
2IOwhwrivHvtM2QqG2cBbeIeIxo0ESLVeo4lLzLkBfX1Fg48bS4bjDNKblC3L+Xq
qxPiK7g/OVsJwpqZi1/2/gLVYTdBMea5ZObM5LKEoIB6N8nUfkHPycZIsvFpprr9
dpapJnfb6T+Giwv1M3lxsiVWdyegy9tiXmrrVlc3Dd15O+VNLWU5Lryvc6AdJhWz
BWXrQinrYvG0LKzNrQeRCDJFQy4/ztmJlb0/MKHlRVprwoI8rH2ryrDsKuHUoejc
mCVX7oItYI8m5QZRDwhFxQ1mGSps5iN0gOYJ1SondfJlfUAINL/de060+O1kQGY2
9mNPswUwpI0BIl531mXwwwlxoq/fnznHimL1BtCdnN8H0purKkgOfG+HBhQ61XBa
o04pSKrFbMeBvDlUu6EnUljDK4IP5wO8bhZbP5adn1rESQxExQEb+LdVKVF4mLdf
f034GQgswYevKmDXt0QbmGfQesCadOuwmmzT0I115ipIkrP1ZTnBq4I36W52PBy8
8wTTD23suv4p8e6AfvffSpRYMAj0SsEYI5Mo7uIXz1jiXnzzw+b0WJle5zsyXv/x
jXrdFhSxYY+ptggEA8rWrV5ranKS+EyzmArHghICRkui0+9oMJHDwZmOj08IfDTj
n8OYO97ZIqIOJ2UakqdNVxtE7+bTCa07cNusl4630t6wEUrfWO6pre0JR5zc/eut
2p/0QCWLR4VL79/J0VMhKgWSmFsc5FnOUqh8805KRpCV/Slbum4WJMROquOho6ru
QDmAjVVP6YsjxzSnRXFyIdItNRnmPFN9sZWtFiHPilcmGdzd+QVadyrPP8XFJ+qC
OpZhcu5+4udz3bT9J4aE3DODb/w11TcW++AOnbbp/437Wev24G6Fv5kM4eLSXGQT
zCdPg6LMQc78N4mvwHO4hEXyXL19Ai3sdkeX9tqm7KP/k7FeQrbwDr9cjeOz4pgW
CcxQFwkptOaBd8k/V53yLHaJg0v7EfIRNn+b5pJUeshpcvh1qQvq48ld61YkeaY5
jeuppt34oiK+2tDp0R0g4LJ3JWBK7a6KqVUNKXeOi7UzC/qIe2bNUbkKZYgMqQdT
FubOe9HJms2It2ujIGbCAwAIWWC7ENRoqEr+J+ckQVpFinsP/4UvmCitvEdYMbhW
aaYz5f8xC3lTCQ5T0MAI3zKGB+YeN0PEnKIYlykIOa2YstOE4zBaA389/f4hvQtK
xu/wizJbO6KYkGjyt+ox1P8wlwkZOOryHEtgkZE15tCj4huY0cKNragvy0IUVo2l
ADtAQeWxccq8vP3MMPS466jsDsuHBXWbJ/t/eI1vUjR1ohMIoQ4EBW9Tecw24M7w
21bwSbEetMF43I+gd2oPF9FvWAo8QajWv4YK3T8tQJVIOkVPFPoPGHt6Thl+em5N
ENA/Movr1+pmQpyq6OThaWBogTieP+hbu1ucGWyOhAebGPYmjfmLwFaYN7uWRz2c
N8TiT3dx+GHK2AHC0ajTJahE1Ie6vym5+UyJatPt4Knpo/BIIBNN4sB4acex573I
Wxg5LNLp594k9AG5G5SrF15I93IN9NXUwkLHDC/lgfmXax34NknPBzXUalTzSo3U
bh4ZNMgVD88n64pE7xJjTmkewwMPsbuKEXkjyt5hybwJ14KtqDYzepg6YIssfoED
KSveoZ4r5JKi6FjCpsCpgnrkCAx1X7uTJ8LHaMJoNIxJmR0IeVH1kJRnH+UcN9r1
EtlTaYNxwkpKWttKs6G7I/Z4RBWeXrWTOPkBxE1Ikk4fVSEPNHvh2akXz4farzsJ
96XbQGIiz/8+m68InOGZ5qyeFarJkl1djLIr8B+k70moXZmDJejUlUQTloDo1DB9
zYrn5zS8A81u4uGawewk8Qij08TFsqMeLty5z+JfxZEe4xuhInU94SWupvNf38KU
mFWWtkvY63XlzU8+2Qu9MQ2NeCnpJwJWwsX5kH1PkIYGrKKYpygXIIPxSFsI6Le8
eAF+oYkko1mlsuw3c2eZraN8rp050ZFlJMzzgWU9tmm9F+7mJDzMvGG5Gv0cTDeE
/hdyLpLAj4uwgiEEt2Z0SkX7Tkw1Xs8fx0Q1hioe1NIpzbPG5TZqMDgfIdLLeODz
cldJBbFSwOQqawIFsZQ9v72QS2vGFNGBGi8Grcnzi4kPnYk+PRhW/cJzcFSctJUz
qpaa0oaFD6nLCRUIQvhl0tO+yM7cjD+IkpfSqy1Y77eCcuneQIzqDzMyr8ys49iV
B67c9Dbvp8ZJdQ/yBBXfo4R6jFvaJqZbGh95hB2pTyyV10/GKSdVJgGvEl36wmzx
tXZKx2BjEgFczGI5fEAkzy+T23zhT4RrI2BsxkOxZCRBDxv0+WDBSnDTZYd70340
4YZwKIOReOO5hSAITymSc387cU6e5U60VAb7xnDUNUd4hY7oxuhy6gtTV1G+W5DN
JU764mVrHUjHisdLOb4RsmLauEdgoi7mw8jz9sAOW8Yc3jy9gYo7hT5wdWDF1wXl
FnWXnk3LDYqsUL48Ta85/vjTR5o5amQ7Nu6KcUm+lXF8cndIWIxzr+ROhFL6cpfO
Z3FSUMLl58vd1kQIgiNz7K9a7czjJC2sdSVO/eDcXUIPiwn32Mv3c1ZMOctXiEiM
tG8lwNKsGJ+3XiNMAN9wmWClNcgTV8Kc23UkQAlHsWam0km5lI0X4OGEuKB3sNSU
XzcfgvEg+Yugr9mrN3zh3VUCxlvTrd5nge2VcLU4DomAHP8c7rLMuIhUNlw16I0q
ENyh5pMtA+a+m7VYyIQvvtSOV5e9HhuppQ6Th3sgl/7RpHW61SDOld6wK2UDM9El
FyW+qNz9qKLMOwxx94DKkfs6unMmxZ1a8px3BU7e8Q/c8ohx1QCKgpLX5bUasA8C
Pv0VE6DglvI6vXlBg5g17wxYEEUpftwp/WfkSKIRWB6vcuxy5zpcpejOgyjGiXyd
8riB3fJs239ASwkpFEOXevE3NB2ZZonyzU2cbeJuFjmPVHkqIpjloljmrrR2NEUp
ra+Cowm+JbY17TqJVI4+7Ciwvirdg/CoJS1aSDtgbMRM2mkt+JQMpIkUoRifwy0o
4UapWLBu0jhJDvADiLVDIVxnKH2LAunmDknQkYQtviaTiES7GdoCnRHe/ohulBLe
MH4flh4US9o6vnKE90aug+8z+hFJ0MRSY3MTlw3+XUMTRa83G/Ss3w99JfcGggUr
dcsMiGrjQG2Gx42No2xkUg/GXa1GWFB1awNUpxkwRAzGBUaEjze9Fh739u4utCFX
pduCJfKahqVPa4NGo1vmOgLPRMkLZa1jZackQN2gPDsEc3UMkTjF4p3xnsaljVKN
mCPRmEAECYfd9l/H0ZC7TFdtIfAEGpd5zXPYZcPAEVNmb0n5devWKv0l6/LRENhq
e7dNgoka+XX2LCuylhQL0Y8i1nHcKTPMlVaOtCiKuPtTCcNuOvoFmnIvPs5JV5NQ
LgkWwMv3C0FkgH9vzCMjBXBDDuvDlDnkU8wF0PLS8XiFvRzaZGEBhugfaQ0drVMw
HF+md0J28v7D5qsCDe0+ma3fmEt4mgtjwz79wxa6gtTMpxr2k5Q5a/76CDHdrIQD
BX9Sh23F9Vx3ukACxKXjAow9FeymCVI3sejP6pFoPHSnuiYYYRXPDW3vG50drQkZ
XzG3HGOCAmZ8SKw15hmWyZ6YhkxP1yBF4Wd6LUHZrjIiEkBeW1+wArNFTxU6BS0G
rOirfkCbkPMfPv5jHAfXfygZLuVlnnvt77TS+0d9cJGvr6QxII14YvlJ0NgYc6E6
cyynp18TQW0cpcZcFpQNO9K+sR3786y1qwNQc/D4ArcSIKhB9SDBgIDWDw/AxBxh
a+9CG1ynwk0y4VhcKzWKbc+fKPAdsJXiXwUrz3CJPMw7eECCCCazsEemY6g22f6C
HyU6U9fvxEY9J/rQ3TCvEBkRYBtqIUVKN4S69EZwoxa2mblEh3Ahb1eguFMzaBQh
pTkzKq57ZVTohTiqIkBBMh/sUHbG3NkO7q5KxNRBarh90L7bTF2PpEXrBsA/HR47
ghZbJrbbiexh4fREdxyfQWtq/CWX5quK8I+Gc5DXVC2x7aBqrujGgMwgXzkTQ6hm
BhfnX/wWsGMYC9CaGqMOGoP6FlkQU3iA/5aDgwLlGWk4Pv2E2olpiW0Q0qp2iWkk
7dM5TP8Pn9EqZ0b7kLWKMZKU6o+qdvtPUdsclXLsMviolH86mvFOdpAH5AlQAF2z
fyVRe74v3G4YCuIjvuc8APk09aKykCtZIIOknWk1OVldICrOJUI2YOEsuJ7YgxrY
bFsdU2/Dzxy0ldZQARJLe7tI/QgRhCN9ctiCqRUDBsi5+KYvu2AOTMa/AlqF3WvF
h/zF9iy/zP8qX02cmjRpX52r959EAx3g/D0AL1KwBLwpCaCwp+Mikve5QzRFbaU7
b9BXQrxMgSkjmeRNGOMdNMRGxE2kHUO9w9WbPjiOtpWyNVlL041YVKuz1MTWz38o
4n37SJuzSWx2WlPB9mtJy1nrpmpPTamNwK+Kl4FADMGX1MAMZjUBJpqzK+8qiZt0
cguXjzcBItPLkMcyREhbY7HFGFajfoBg+LxaX+BCQl/3fMiiqMlPMOZdXr33p4zI
fzC16tY/lYloz99r7gZZFLj65qBCxA3m/drT8E96/MfV9cyQDp1ileAH0WtReW28
tZ7KxlTFHaZoeTiPFW/3CvE0qN1idlqdXtbHcnGn5E3cvtN0wTrGd4f94Njth2jM
rz9DRqneD7MCieUKCkMoMDz3/F0/RwG/sjVpbBiWJnRLOUXmE1/bj6noxGyG28DK
nEdE48+oV0qyQU62YuKsCmSxyfHqy3cVGbhkZktOh+qHXyv+Tqe709fKOQ7kYkhp
SwI06pXYIAsN3uNS8ubEINWH5XIT3/zA2q1RpGp/A4y5GfYrVtdjdL45guSM+HO6
KgHy6uSQBKCnO483DHrLnOSforEhH9YzlbhjZ1PSk/KebxgnuHE7K6mxPaDJILg6
qMmFynT1qos58bZQvQl285f67D0IJSKkHR6aB/+ELfSB34hVLTswIH7XMt7SfqbC
5BcEJeg9mLhRJcYcYGuWIe/R5BvFo5DLBLepcuhJF/++VNf+NakNEBLx+6GlQQmq
yD+Ks6rrGhIztxv5DKlXDerr1ZnUK/DaloRX7TcYsJsYvfPQ+BLT1NXA3SDlShtD
uc8EtRLAL0Hq9iLgNtl2oPyfVfHWqQSsP0fYrKV6pDG9g12qfnvs023gR8hAddfe
CAuNwN0O5ipWHaa5Lopm2Dz/Zj5NKwPbS1om4QOy72le6wjbtZrIUZU5Y0ZYy6R7
DXKZbSCVnUqz/AW4cZT8Gvt7pFHAwLEiflVrbZrMMDHjZzCfAr/ClXp/iWRbWzHM
+KtevhzuPy9ya50sLnOOSW8CJv3siY23yaQm4xb8M3sHWkDYLKcVV33Gmn8OVcnn
yCpaq0ixdbRIaIgUeV7HuGcmsGOc0n52vto5O4HsoyoxZZK/I62I8MiEm0qgW0mF
mSrsljJg+41oi6kBXkPOd3gv9ni1ibNHMx5PRySSyRu2MhRavJPnmdZIHZ2Bc7GX
/Xwk06ypu7ifUXlRaBml8QpdNenDIUEdrwpAedr9yGhifO0i/DYDSBZKI7GB2xCv
VrhW0y2N+kzilbHz2vVdeasfjQSuB7NDfa0S0dLOrrkpePFSg7Qf+qOnSToRSDfe
pgoUaeHdmIh3wwY6gm4+bvRvkJ3wDato/Pn5d+FQe3IzR7fHEDPEwyPx8HJYYfIC
5b4aB75pny641ReCOdlK0sirKVpOtEVsgfXCGgdajz8VPhlPpypxa6ShNZQ38N8L
MqLo5crK4wttdYPWYkIttNNr7XciQC0LaFlZgJb5YRiWH1oNWEz+UeeWu1onZTOc
uz4ngjpIdMb11oBe6OUm4u9HQcdTNYKk6U0YsgISbbVmptT5mbr05BuMGs0dqTeO
hcp3C9xrz3NWuNyIzKIN5W0Pw3hVvgzO4Pz9uV181r6eSrhkCOReuSbsGIGhChcA
Res83007ANpipvk372INWtD0h9DnwrMSlILcYEzpSUo1gVLjkdyr27QO6cq0SXi2
eTsL8G5AlvOXqmvLUvbOKjFWgshAHbcHFjQBxb1RVzRtdQ0W55XE5qkWoQLM/3I3
//Zi4bX1op3noyXffRI7dpg55EcRlXGbkOaqQO8sQJSvKNie9NWGHPg6a5P1YR9D
VzbbaHfmC/4rHy2PO1TXKbhtxDVoN3//CaodncKeTkwvhM4o0HhZVFh2gH7Lt3KW
8zGzuAwDdAlcxVEL9kBFlncpgTSZG0Fa/S/W/fT5/Y9BKqXiNb66W70hkLHdrby2
G+6UxW0AGDLxTKpoyUbGnHFgQmCALRnnxBXMBWRKrl+GF8plr3MuuF+N/0Dd9ngD
7XjTmRMX9o0sKUu/3v/yWP8pxsM3kjvKfKf0QsX/vXWLv8poo8SWQ2tJKamOgHFD
oKyB8w9/Pyw/MfAKABC9XmNC9v67W9AjjlUhkonSm7DD2VShodN9IGk4tK8dWQ6d
87neh2Dz6rWMk7vk8S8ogVfDh+JmVPROqTfpmTd7FlBSTwwbzl4CfkXICbO4AfZ0
Fj/u/xEKOcD7d9Me8M7Da6Kp9xYaUptOmg4deAeScgPBwyJDwwZ1hlt2WSHlfiuO
GHJz9YEnWLgWUv9MLAZApnZvOshRYXdGwsHPNH3U6EIiCRcOWoSXx6CzMOCW73Ug
NKjE/ZwMbCw/CjfZl2krdFkUYRg4ocK7x3nQVdPrR5L7h6jI5GcfdGbW4kXWAid7
FgyKsCfVV5HgXIHJwgM/0KoC8byzubs/2kTk8y60Ec0SScnIIxwzGRbkpPzUikCy
NwsJxokeezqxtHbeWt5Yfl8wjpVmVjD2jdCrZ45nEYEdsyyCuyLYaJCE4wG9Hmbh
+EceFZb0WE+rhKAahFRT/JO6IHVvwCcjpp1xWalBMy9ZyBbhc6D0EYLXzxKJL+kA
wd71aMlRWpeazmeRU0BLUZvXnAm8WFe1ION1JR5voOIzUONtyL0jaouJGdY97tGH
m3UuPpvRUInJaCQZu0+LGQ8ZeEJs0YVT4JZyh+Lh5ZVo5wzeHfk+YSBtALx0niv9
6ovyQOIrDR1VvExVWXtNWcdcXDWAEr6e8HRlpisDniSzWo0z/jPrtHPIlWnJSIC7
Yl2ei2JEWlCP3XFwUYmDDY3RWR5Ifx204eKfnZBU2AiGWKISNqM9IAH61tqxMqvl
erykcyOyOfFq6Rnxa05UnvIczcb0b1YzK966JesYx7ofl6JB4gdJtI2O1eMRwleF
qGrAPp6rQdkFV5yuHe/6EA2Rl7JJWAn+5aqeEw+0bKK9F+ZmzVLTvwAH38N1vjhm
QfT8NsKLzUwRgbdOlCfCakvyJOT4wPVxNIn1nNsvpyj0TxVtRWbkmvLsVC2idkEQ
zBBTCwSyksNnkyyocdalQB9yaiCOVl1eX1pc95/0fPIiFf8vpfQDdSc5FQNS7p6n
0L4Gz+bFCiQMfydPlJkjSbI0AC7vNtW+yB3vIcvHOPGw6fO8hLPB+Lg0ssULV6ty
k68lnUxRdA5Tn+G53UOohT7od5MVbYd+mQUxv7POTJJ+BU7Uxw4K7Khy5Jc48iYE
NDdTf4nfgZTY0JRDGo5CMZoUA5S7yin+h8iR8bwZ7g7DBkiRUXaRu66/S7ay/4r8
YNf/WcbiT0ekWQ60ykZLZvX0wmRvMZ2fknGsWgdzrcXk2izf1vrIPO+aJ+klhFKo
E2qeNTpgeAzDiLHL13UUyYfQ051tmYwot+opnebgCoMwd7dT7z00Qcp2RYMh3lU6
lDfyFiIdqC2KgNzDehyH9dhG5mFSEhIwlObRvAlbC8c0vPCE4TheVJxmZWXgxyzK
zF93BiLq2VC5gY5KvG1kHIgeSWaeSpJCMpboZs9fEdbSZ6U3H3NAhubfC00mU42/
QDbs/aWsMUJtCszZSRqtZBKcaLTmQryVMPK5TA/vD1l07Pn/OYGxQbfCVEzJLn61
VoqACL2AY/9k537edJNbTmbElk26ABdJT7nzi3mEuujKhwzdAutO5Y1QOsNOF0AP
j2UR5T+17xvV270tMbqJP/ib+PSgT0zbnOtbzAUCul4cv9stoM5YF9ewCAb1azn7
/qCPxCoL8m9GhSvPFawhzhmQMkICwMu8G62QlIByD0m7L0C6G2nJGwR1qBl5aMau
HQdhPyTAqg+2UBlUfmvbR+Oxp0TmjzYJ86qu2P8fAhfsuDjvhWqbNQAsZ8qbikK3
NYuIqUpAw5vAX7tIINgWh9CopxvYfHUoayEjJWzYW+Zts0ByY4KO7FOFYuSJMZH+
qAYXW42Mtx+7pKlj3i5YLNFwm7Wjs75IqEUmRWbtsJuPO633Za1f0q7JG/Tu9Qw8
CIoka8LDFV7Dnkf0VledQHbrXCJ8gu9zUtwp2iE5vRBiS0CdpxCX9ZMkXSN+EWqo
4jr9tlQN65B7PzFpiqlx6emPFz0mTbEnoZ/rptHQilMOGghI6FfoYFniRLva+70o
JipzT79D8NbwZ6o/sm32ZLENS/H98/Xm+WXDu/JzMfpAjvTweUMAZY2enF8AG6NE
bncn6nQut0Qtr77wHmdeQRpUdvIP4uPeKqPJmXrdueqd/NYsZjWgckIuR6fqw3FJ
HXAnvEchIKkiqrNoizKLory7qUvHJmZr9NqwYvW4K+22FbS+EC2NDtZLeUsucIzW
pTqDV92/M2k+MbvJFFTLYKPPX4Z/3e2kDGDFiS4raq11l4oFJfu2d3gE/y52P5oB
VyR/Gmzem5Ve6ApIx2cW4mZSLdGCReR0b6rbgTwyhn2qoO0ULJtmS7wpBGlZYv7I
8qgFXgeI0Ynba3HCjgY6RwZTROGjTfwoId+B8GFpvNo91I6ZqfERNNZO7JbUzRkc
Wedj/mgXSIpAIO9mb8WAU041mn5lLHW0xFPRge632ydny+22l/Xn9dt8gxd0jN1X
P31zrLaY0PSGsUp8G+NpR6ZTCN3wdhVjFVu1Jif9MhgnB5B7poQbZGtarsA0LV5C
FWpqzJ69IciIeLG0NSdx4ZIGZ4gzTYgaQ53hQy7r1D+a/ThtBHdfE2noWRiwBIVe
qezIcqZtjXzeXN7UWA9kVUrKGf7FGCDhRqA/NySapLy4KwsCQQOHBO3zLyqgj1AI
3UZb7vSxpoDeS35GewSBdh4k2Vg/SplfDn8NDD8hSnwNVsWIAu9IM2dZiQ2mYpiW
D3qONtOV/Slod1D8P0kwQcib1q06EZRO3o6WS1oFQfWpqijziNpr982aZZ+LiKP3
O9IEyHfqdjqjevFvcjhwO0/2xnkWVphIjb1/cI3XYIro78M50A5XA1aTtgeuEiaL
xaeoBtkFTfnL//uWeUMt0KeSsyh9E0KiWNqYWWaOkUGSBOVbd1s2q6ps2XLvuPyy
sYZrrVP3BjXKaZj14fZSaJgzi+eSidM4/qyxQkYhchDZrjk4gKsihyDEGqbAQzUc
YsznYK3xLcokRCtZoxVkuZnI+6tDfkzTauMK7cdY+yai3rQ9SuH6DzXWfViq5xO/
vL5G689vJlKdh0tmJtx9m7NVQnSvJqchg/ahqxqN40fePt8HLWjQgFRwGvY5Unxk
L6GRjjKYURqoBrerk8+G1sMQpgMMfExS+tcQpvL9ZV8RFiBXFe/qiVKwR+jOOOtj
/PQkYxvTXp/8Rwya89LRRxaMEdg3UIDZ7eu3D6b4vDZj2lTDZHA1WPXgWVJZvqrK
hvzUthL7jnN1iaUEvSFfeDrr6Tk1a9C98zLFx2yCdYE10M3T9V/aNUP5LkGaH4hI
7sPrYV7Gs0vDO15VrZ/XaCOVqyEF0KjcqlEf/qCHGEMmKsris886vvO/4nijCxDt
6FuksTvllIo+U03kKhC0ymsrqFV8dw3QeGj/X5IMqzjNwa5sAigGIijZOUVxYjhS
+mFobTQ2mjpAOPerOfWI2RnPZR7bTrqK2YumcNw+v2aFit2+3Mw1qurbAAQf6Dus
iOlUVEI3o2iG9eLGRQ5CJrdM7jE9Uyj+Rv5E6VEGnZ0Eg8MfltoppNzKUKz7dGKm
EJw6cCy3X0w5XRdBC7VR5g6/EUAof8vfB7NxsVfLHgoUHI8jd+JBwK2JmmX0SIci
AloSG2pLwIWKUN/FZRJsJbpag6TuAZuzSzh+eUefFGeOdnCSuF+dIvA2wbOjhhMe
r+U8KLZlkKt5hGXERwmm5ai2AoWhfqIidTn1BvNpqxal1P8ErRiYSV8OorBe3WFv
gZFVfxidwBi1vh6DE0en6iDU3xr3H/F/skHVq186pV+mkOLCcyzRWM9ke/JnZPT9
exM24i4dbZ2OvB24033W1lXcDJLjp4oE8veODoG96xW55YFk0WGkAVg3WaJkGOdl
Ccr9W7PTSAqdLsBNQ2IrJKYHA+UTwl3IVr4l+8CiOtdQiGs89qJ7TTWsQbifLEsU
t53PbGJ2jy93si/OiirmQqBpkLoLmCGgRvdfELXUVQpbREIFNo3AywVApHTvlk5W
GHok2oOFVU+sHw2s6Jhy6tq44NFPXlQ1n5eA/ctJlIrFaoJN7NsTORVg0QmHiHIV
0QaLw+aKas6CQ81TC5cDryd9wyCoX2GCcxhBB27KjROvpi6OuYidVRgxVWcPJRBP
gZeADPnI397VRgUZnyo9JAXC5leCneDO8sDEXJUs09sYhzzCXeniVDy9fwXec3ZZ
2HFlYEaFJRbAUaQf5Ek0W1n7qbrv6wpktEmoH3CmtOk1PZEBnSHaafNSco4rblSe
PjBfzFxll5jxpqaVFDpBxSzipbHZDIowoHgnkDaRWrPf5m4viFEnlNG8oeIQ5BUP
qspg9Ryu7sBl5VxAwWDNjzGNFFNZq6jjsHeqxZ9E2I2yW7XPjc0qaIC6NCvCf3xh
qPFaKNFUrq/2V8kRaKL9Nnxa4eoF8fgxu3NtbTOk4vXOu+YPznn0BGNJKKEFu5Lj
QmtSYge6RVS/N/V56Ess7YrSHLN6wPUtgBugakk+xHREAeZhICQZz04nQcOTw7vG
SxAWvGH6oQddb/mZCq4A91fmoZAEs98tiaFh0zx66rOKC+K9a66RhqLP0smUvO92
zEBIzEcjWyCVD+o0YPihZ5dOrow8E52LM40T/8ybB9UDQG9cyVPRYvRnWxDPOsCt
jEv3F/cZa76Ze27biPFMgRMJ7pV8QohftgHzEU9OTCNZ2PjmTxrLwbhEvwLQBbgp
z9/WsiW1mhph+ozFj8+AU1VTuCtDFKcn57mIEkJBsFLTyiR0OjD7CF9bXqmTrTEw
kYZVPQeO49zoErEcLKvH2lSZsObvXmuEnJlOEbSoL6jaOLlqJYwUg+IsBRwxDLa/
Br6rvBrNGLo/xRGiFD6ocvsYai+4IBRdwH9nueHxgnWcyKj5nbfQWztSVIf4Po4L
SjInRTwlBWmZH3dbst+e6S63ehMp6SQ+aIuvNQlXEa7pM0vO2gcMrBoKAlP7hiFh
b/21evDLpv65pj6Dw6u4ZQrvivb6sNy4WOLjMTscMVXUTfNi7Bk2PHn2X/1xq4M+
gaGE6tb5yJTVcy69PZmb1A6AkECVWIYzdLdz/XE6X+hdoHM8vUsdc07XPsvImD4V
t0j5RI6E6OK9I4AlhHSfEA2mY7CGsZCziKsVLICDnCwa53kzdfN+Ep/gbmn6TeJh
4AaPPZ73uhCYi4+3h0KV5dXhebQ0cI7zGG4GAqd6YA+24EPjeEL7RQBPzvgFwWAb
w5n6nRBzob9n1GKpggpPlm+PAziz0xu6dBanTljcMK8DmwsJOy6jf3mhuDYXQBee
KCi7O3t8CQIGWdCmCAfYkhxjuerOfU91DCv5jmjhJh0taFFO4puQLaIZqOLl3tPq
sVI4ltuAt+a3FAFe+bzqzaO5fAV807UjaFrVLWPwGKw5NzVZmUkZZ9/KS5IVK/YU
QNXefyJ5arFxZCYwKrtv+1/yHoj5Ucooipjr2JyRb6Qo/m/q5gvjjALN2Q2oJsHF
gg5hm5cMm3C/NqVsn6FvM+cKerQozVo3duuU66REwQ4YnecMGDHgExS44LO56R29
fAZgInzp85Qba4sAzLeOYhMHrse+CvEjrzub5fxa2prRuiiTvBjZAhEwjQT2b+y6
F+g860Svkx8x9TNXz54jVeDwhcYKa0MZl9wKO6eC+UvgJqW46Pk6gY4la1gZdPeH
p8kLTaaxtSupX7609V5Ovy8y4K20R7iyxi116fmoutbCJBauakFVyEeBzsj7PtPy
tzdnGfG6K1WxgpmdESda/KJ0P4wlw/QzcLvivjv+A20/nzi8lB42x97i9ETxjsry
oW3L2LyV5c/Ll10hnbxnj8w6PYD71PBA+EtdAIh4o4QFds5ysFCzbk0ZbzzTB7ok
rjwTzgy1dX3e8gPSid04aGt40TkfIQJGkFXcU5ODKLmY/MkGute78tdyPSeLCC7y
Ixyy0BtlP89D2bgnJ9omLx3S68eUTxvpW2uMoYKK4PSLAeA24NXoLmL50u02nva3
V7K9MLnOsMucZQTE0l88Nik1EqBsDIddLDgJ7qKgPg4u+mdzsGKz3SEndwerM7qf
iEvGdK5geC+0LsZFaXHDSYmfedgNWZLFTphc23S4H9DfW1SuImeoQb8Dv+1g9K5z
sS4X7+zY+8TRn7H3/1RibopcsDjrGt7Ifgsqr6oZsquEiguk22cztRZ7MfvYTgD6
egX2U35xsZa/luCPQhVwZckAKSvrGduK2etuxbex4y4nf/qNZRVETDWeEAS8MSo3
hFcTuKCTKq4JJLo17qWjZczDyPR2GFF1sYIIUiva8lZONg2/vwLbqGOOfO9lLuMo
6NrRvqi3x++gNcCt8wFMjRZ4Y/Acj2m32QzLLqRbOGWShPIsZddUL4d+YxBVPd86
0mQAWjuOICpM/smPxYDvR/WGmY9WkrcaUGRNubf1xK2Nm8D3FleQ6pJDRyiVL9IX
c6kW9MCjdY67xl4pHRQUMhqIH8zPo93QTHL1VxEaJcW/itEkHQ0JTBNHjXcSH6Wn
pvjs4uNmmHoL0c6i96GpN9o5kUsa21IFR6tYDllm1BbXDNqDZ/wFUl285oTS8F1N
QANhjw/btUhOl8Htg4fFV+wpfxzJdM5WU/I6raH21L+6PZtNYG6x1j2PaqnnkTFa
ZV+4mP77eXYSAyavXauKb3cH9FvaU+TOYE/uAnf6J/IiJOtOvK5vF2F/PkCJRhx8
zL925asaTuAeVFoBvU2fhXMm58MP60vwd3MksLEYxGyiHPTaPdUF26OPbam4jFZT
SGZ97mEsYkqyHWbYDz16aIkxnTRl6RFHBXrWfm0h90SjxLlqrtJJtHBm3/pw36dm
GuZhv2WtnYGfdJY6y26bOz2djK4C2Yrl4nRBZ4sO1tghZk8o9LwHoVvowenC8CX1
OJlDABboyykwJpITYVjxZ5NRSKp3HnyjISejExKFMB37ZqbLCPlGJtfnv0FTbG1l
O6LIhgWQnV7Q6WJsHZ0rz/lueIRincLVzZVmD3QM2WbwIs5oLOha9g0qAe/4JfIU
wAyWGSoQa82u3P+haRcg+LOia2RRL4SPNDoqfJosH0j50SivFAjZ8O6xPLWDEhx5
PUXo7ND6WVdOSdVM1K052ml1V0i+7p+P4deDxl/Ojxqvj3dUNScfF3gXWitVI6+m
cb0OAG9LEADRO9f2FAId/fn02fVuJXtSXKCSzd06A1kHZfpv9Inh4dRF0+AgPJC1
PasqHPKThlk5s0QS+jP0pA9cMv7lq4tVnKLXkqSIthlOotlvdSkicVHqzL5Jx9ej
j5sqw1cwbyDIHfnUChYMkSN36jHAsayhTcUMcIGOd6u226mCIoB5c60poycvh0Mh
YJDyxhHOtlYgkuy7nlp2wCwjhcYIGDBgOcJRKrwib3cc7r96miu/QaSuzzTWkSa3
36t+eHjN72grgb9qEipT4mzHg43+5xDFgVFammyRevLq9H19tM0l01WZl8+vnu+a
vrEDxTTtgc7M7ovcKQMmRFCj6aGcg6jOj8IkltczT7u65WJioL1UTDpoWpzbQZz8
mcVRoUZZSDNAOZanPuSZd1tS9rZXJtoP3hdslObOr2gFUCSnjEZf3PY4aKoBGd/g
zfjrmT2d00uS6TLoVmAARIjyK1mfPKcQx0fsgSW0ghoB+k9BhsTn7yBziON2Pmy3
DrFTsFb5WMfJ2dE3UOFu2qZDcw1bDC4p4EGfVbah9UoY6688T2AhygFpTlPLxiyz
951dUOSz0fVSG6ggBT50zHSDfgKTmU7ELmYb+hz4wD6qAZy0PWuoCH3NmIYk2XA0
fayDyi7HDV4j48D3/ekXBoUPEcrORB64wRcH9c2Gj2rc50DC825fo80WDEwayaYo
mJG9FFDAJrJYFp/br6re40tj9tkXKcy1jhLidwcko+NofvtviXAMDmWyN6qCegc5
cnHovIbICJ8GU/YIabpwzmnub0rsArKiuoBLE+SrfzZlrgZpvWbNLQ5OSk88rjMX
P3zRZrJzSivtvTQ/yZdq2+pwvbe+iJlYhxAU8KrJTFSyjGF3IRd/NDkRaNjeBdOj
f+bRVah+WhHGFg/MBOjQlN+2TjyGXMLOA0m7GrU4GjFpVf1hkA1S9wSno3Gslv3e
wVvYeSKy22b73Jjoqh+bU7adxnANZB5J9X5+SsvWpEJA3zTX7rDS3v6YSzWCgKwI
kQ3n2vJOzYp0VXRZtFxwhVMpV+cutNJbhpYB+2OjmIU9x2zH0TvzZnRT12VCkjwc
0j07hlGzXoxIsYQPqivnijf0C0z6nYIr7vpoGGHQl7YY9J2V3u6csEKPzErLnPSn
F8TalaYVfKAVBBjvsNHSDKzP2pS7eedfgxRpECb+hBpqrpKuXjX5PgYOQvKXWZjN
ka+42oyutBlrt+9H04ZwSKSU2jaW9ZNXLarQhXRHyYs5Jy8PUbm+XVllOpMRz0gc
gz106Zw2FfDL3IIz1kfKheimPohaLfH2mpG8ea5qBMgdES/g97G56iLSxznLd4Bf
9bPdgsH2c1Jn+USTCtZPg8JAAvTPsRwN016Ac7SDrpymVv1a1VczpE46opJj4FAs
Tbu7Tubsj/zKDO/19jCSKFlVf2/fiTLNmkKdeK4g9KgMR2FpLgLvU068FnTHU4yb
7v1KBwtGrBiCnO4CiZmr9fUcGYmvvxCbrOh/paofLHJX/lVVfj5awUoTbZON7Wzy
ac+7Ptalc2jXqqVzTe0dioDz3rJx6o6G+malpYF3+1d926zXahlWDpptMZ6UF1Ey
bN8PayoNwtPzkxx/bv42/sseXJ5g6LA1x6iyjeN+BAHFiF6EudwAtC6thiHIgeaA
hii1BSimk/cRrbntphTzJpNAnQArzxQcFVFvMJcuIvGZg04wDNx0T9tNtHzsOGX7
GQfTjHuvHV9+p9uF7HV9gCTJclIOtCVOQrciOU4t4e3tmr/jmrDwSYIQ67tyQGfL
r6oVxGMXglDRctv5hscHzk0GXFh85QKLSbsvQUus7AmetLfvBPrVhqpsks35xWE9
Hu9W9z1KFy+PeZQfIsG9d39Jmm44YQ8ROfeNPjNQK8fdKVx+sf7S+A6tKxVvA5e+
rOk/vHIj6Gojc58a+8reIezbBakacMyEh7HaKWCQht+QJQo0CfPI80JAhrTfXCtg
lymM5JCIgMl7BukVfD5/+SFbyIlHEE6ooUrIJCCuX7/bPSRDcvQbTMg0MGmbGOMW
FDM14xL5SF8F1xHYye4IyOjNRevxD8SGPuzCQmNlDe1zF6MUjbv27RhgjV/eAkvs
miX9MK3h3BA1PMSiXkE6JKI4bc0G/hW3xlVMu8GBV1tfjG8MexGANZFpOIAjvt3p
09EG70oVlTveRLNH0OYyJZtKCW9Wfomltd9LufH6SisSfaw29CqiL1E+0dlD2QpZ
R8MMJJlPdAoZD4J63NnDVASMKfJG6WqTMFAuJmHyAItDvRek8xZnBDMXnf7uoPtm
kyGvrggLNXK0gMXFgRSl7jh3Ygc/ipAdBm47XnJUQK7Hl3mW2Xw9YEb5k2DClRFI
XibkLDHxPy+A8pLYXbd6wCRFLG5dhBe3AsDMl5iS1VYWtv6Ckyjhk8wM+qpAKKqC
4QYBqrYPX0Vd9IOUfxCP0/cI/YsVSi9dpj0+l4IHDcpua2etrrkrgj9O9BrIBkGY
8vdH0VAodXssDutRBD3/6AQqMujO3qcb7zLF7okAu7S4qse6rg0LeFL6dJ17LkQQ
HzpV0kwFpJaWi6kCpxi1+tuvfKTMqiLpfme7PjqdAxrycmewd6JhvGBpwJmbKMVB
ISG3Ele+PEbzvVZxP6/UUzdBfTSjoQo37yG0L2KKkLyqTyTuTZuapVBqnRG5P1XG
amcHExPgJcunNUdjKSlbvoo/fLKmWL3VnxWi2jeZqTbk1vQFWBHCb8ka0UlK/7hd
wRhSQdPDDhhwLnooWkYz1AMhEhDmPCeJVWj+6AaohzhGUZfN5s0h8QXKuKDTyMq8
XdT/Qz1sZoRe1SFB59GbM431d+nSca/d6GeO+Gw7XSzMSp2gGfYnVG3OFN8kHV0J
r9KgYI81hIx8T+FLaLX6XdfqI1Qwq5KV23/w1f+jZH+AnljYntxtHJi6py9fXgMt
P2Y/A3GjUeCbIC/LsViBl0VjwxBXe5e5eZtwouPPPV9eqpVrBit3SoScCGcWwCQ5
dzLNPMVsggzn5+uywk3vtfzlelpAGTECgElDM1wPbSUfO7CFoQCYlDpurFtKHnFo
RGL5XWWv5eid7Y19SuJDUfpPSYJTEkIPs7x3aHkMpzvjMn2BanaI+uAA2EI1h/IL
4SkfB6qJDAP50Y46Y0pW2NhAMLE9RNOYXFa/keozovL6y6K3OvNcn6BsPYWpzIzV
Zq27rq/T5eoyCPay9BKJiDGTXT0rjdmGuEpt28iLUZNGpxdvEEcz8SDvOIs65z/x
rCWUtHnG5ky0IMzzRe27YCgaHHft3xAlyWFQcZoJsPVshWBvYqsBolmorw1GwbGT
0WjachzVxB6FK4YvVIV07/oW95V215G55iwvtqRFWY9aUQ4pYpLCY84bo0V3frRk
buw0FvR8Yxji6ETED1pkN9/hy1Yyg9Ewhz1hkbS1liotOF1TadsdOSFZlEOAH4aw
ROIHLpaBXU1inB25OVgrVMIxLb75q3bJsYj2BE4gD3Zpk+FuhMmqlBAeDoXXfLOl
qdDlVY8sKdLnFIJf1cH2gB/cjF18xHRCxqao93Nzt6pn9+69mM4MYlsmY8HvrwN1
mXo4W50Y753ikzV+cVzyo4QbbWpfJsKZU1FQGvLPOW3EIB6Zk+N5B9VQALG/Aq9y
cCFZERwmV07gKsuLXr6hPqXQabia9XsAqKvtT2/6FZz3oZ7cy75CNiLzbHQ8N8j7
KwHZFaOinCuD9NIoNV62+ZylXO8d2g9yMfdgkSxrbP+IF6R301lyH4QHoyk4KOl5
AvqburREpZNwmXtI+9117TYY54V/xCzlQDDZpN3EXW4oIGnayFSDMxEq45NIFFL0
qyoG+UjuuoOuBudb5jvJ9Jy6MNUYXXReDRX1MK7ZdYVGdMn14C4h6RoooqLuRcfh
TeYovaFXkuvuVCIr6xLZhoqEk7jKgm4azMkZaqY9oIzaaNhEfgNxoMuNeO7hWAZB
6virJd17F2Ri6Jg2C8+6imCRYxhEFZIHLeuOrPnmQpEksVGNb8mS1ik2oOYLNNQV
qVIfeWgsSdcEsWDR5WaMQcRXukpON2ysC+MUH/VDPCsiP51X4eII49EBmJUDZL1V
rlY5RPfGZnIL2tcFXA64wb8i2U+9EKwlnyUZWRMTsFb/TIIiGk98kpVmoThkKg97
1r47/fyxxIN7JQrOCxjA1G51gitpgxwgcc+PMu/CX0I9RWxnaxJPNxCoBhJCGQ0f
ofTK+L+GhQ+KAB90bTpRglOchJkunL44Nby2i8ooPWR17f/TtKvWV96kQ4CIFQev
mRyCivooVn0ionj1eXbfP+o1cV/3lWDeDqvWkrSL+vfiAGNL72o0vSzPQ55lGUuy
3m2LtPxIE4DYtJY1YFiCi2Mi2A5QVOHYXqOCFISB3VpxA0gZGNOeJ27hbO+ntweY
x7XLEtsK9HHWq7ZZQ8gisq4RJ8nLl+b4Z19PwsPLELfIr692oewJaOZWoVA2kW+A
QUWUgim7iW7jqbBMDeQIUbZKk3gZ1c0fdYlY6z26CXrsdhY5UAaKiE2MYpRsdcM7
ScTKpE6ic/hoDqxhkZNPCEJY0aQ0A468EZeU+lUDbOvuQkPEQd3k+t2rg9esz3XO
fQ8aq7mHlCZRIp57s3RIHhWtp/KWYR6aR57P7oUwpipjAtMwOStAtdO9X4GuROlF
L3fHaSIxQM5nTE6sWwReDNXA7w8C5d3QPg8SszxHvv+tWsD7NI/7USM9uYD05y3M
Eb4XThKXnw/eKSChaD4K87fPWbalLvr445wuOCszyINyq8h7sAOltc0CZUhFbR8J
J/vy5UJqP+dXvZa8aDQTNCSLPxudkUOkdEk+jvw8sb1bhmT1S0cHwTkLnovaI1vH
lmPFXE+NnuM0nfEj7p9wlQXNAuHwxtlB0mE43gCVoNobzRafvSpeHlUwbKCMeh4p
xO9M3zBCf6Gr0nPD+Yc0XOEUm+EZOC36IdPtNwGpo4yeuGkWJ1q2+PNN+QRmRTWO
oBULG/qU7WGBBxMy6heYjBBABN2CcAkvSeuwGb9+8BggUN9dD2gP76oaPBkgTxyR
VihXqV9a9eiUalvESWeUirCBZriHD7m+6yCNhFAJC0dVUtDSzjr+uXGuu6T/gct8
v8Sb10MNYz0b38qn6xKS3k8Hz54Xrqgfjc9xcAaKOJJbqmNqUvWVWg7BWnKHngAO
/Di3KouX6T9EP37p4UcbQ5UnMdXQAAtaJZ6khN8XfIrqJ/6TauWmIolaCPoV9/HL
Yd4+T047Ld80kOef7Sdk5v661Ies7BXnYe8vpe8QL+KwoFl4wBcjDgAVUM86IFnm
y00/s4a4Jvu+GD3CkBhjecDlt/L6GzwiptPVCOoe20kjsJ3+zYkZYDZrgUUFOCsD
RNkA5mv1Eo6Yl2Ap0qFD+9pgEVIAs15SOy6sQkxtdjDc8gZkcZwkp6ajXvHlIa03
+PhJmSEKtKZt4g2LA/VmEg0KufZ+g/8uH8Vz6B8rtWBxe/wwiAjDOlUqiS5wFC/I
kVW/RkaYC6R4lZutGtcHc3llQw/v6jqs0YH7khXxmHBsx0mCmf3Y4McxwgYHpujQ
Y5F545hOgmeSzenHXFAmRdWScVXrEqHFRERKgTA5Z/HiY9+3npmDHZ3RehrtbVpJ
lJQxfEeGbilwXSpQe/VkJc+TsbyD6h/sOn9cUuBSovURjOSHjgvNm5XOY0pQpMmy
bMFbhGKK/dhWLAwRrhJ8ghC693qHBnkv3fstb1Eb3kp8xHoTsRIlj6ZkAcNW5kj0
Bs+bcdWiMxYaLKQT/CgTFgGDI1y+HeVVSLN170BcJtL1l96FNb/qYu+qx04ZDPSl
1eWfQSwmoVtGDT4ldU6W3fq2gw74ndkduyZ0ZaQprnnc7OKcgOEN5J3zRcv14IOT
Tob4vq95mLJmmeM+4pzpasaSLKa37yO8HCKsvmHXb5fDi0fzr8u5OhJGzYnf9FuJ
4SeRHcJZ6rqiZkO33jvPQvVzPQTx8Ku2Slr7ZE9J99HxLnxEHDdGwS0PuDm3S5D3
/g5K3vA1wIXdCmI1xFQ+08RfdbVSdYs+qb1aBpxhXhqHuz0XGn2mT5Lsw3OEAvOw
jY8JfFvNS/GIcHSYJMQswdi7Ep5+mXZT3VZEal5340oW48/s6rW0fc9xFkjj094t
Dp+L6dmSZ24kauHpVC4kZTHgFWDaOGQB1TnhAFEbzWvoz9u6uVZBHLzmTHt36AMt
jeeksdES+Lt9VQJJI9weTe6HN9/93+4sx2dz7FmrSkEaKXCOrcO151UwFcxgsc8z
yL8ZOu5hpQuy7/qMOClmz0Vzvf2U3cK4hcPASlvlJx0EiUCXtxdPWSx3ti4U2Yb4
xBmSKMbBDhdJFXFP5FfVCfWcjIzmdKZdppAWBqSYlfgN7QPiazrCgUbt4x/mMZCx
kVbo8VHPGqGq9TCwY6FAOMHduq/W+/ghy9ApL22CHI0xgYDw2DFW9bxgtyTne5iX
ge1icJ08fIaRxV1PDmHIIcC2duvNob7stPp+vLri5xmi/FoMN3R8xiLk74UVrx06
bi87y7GRj1zFhxoK+cMaZhjgNjEEtk7oJA/I0yXRKbQpQNaBDVya1fOGZix08bSs
z/8z9xeQIA+dWOzALTvBesiQE5kVHtw7/GyeKkH5RRkr5xJXokZQKW4csk4kYpRn
+9Yvpf93S5EF/fepfYmAJtbTX6dK1LDKVgs+H6gfYxD+alg53kPI6IWEaWuhxW6K
bmGcY9XHKSFfvl/DurTIM5fBbzL19I22j/PW+FNjcLd3I2c0uGD08T4Q5xdGV+6m
UcyjhAXabF2Q1yYFv9AGY+IiTsZ2ToaPiHpsz/GH8E8I2t9AYBybCbejJIXbal3P
i0x8j76f/9L9bs75AC4/vjL/tv0KQRbo6LOXngtDpwxP4b2776QYQm3MoH3nu/0y
uyU2RfnzLXTbQxKHcu5t5LTyz8QX/CDHeNze6DPBJ7WJakDYO9wLdtoFbIilaHvt
sv7cTHo7QxPO1XTYMuzAJGjR6ySWQ9JRi5ddua/UGTXZqVydzqVUU4AEyA+uTqhS
Rq3WCIfIC+TZcZBE44MigVzbxwALReIlH2X2UxEd9FjMjxEXfjA9gFGzki/1khWx
/Fc8Z9AxZS2uobKHXsRGNhpI0gQfnW2FDeJa+8uQ/BFlU85bRWMVLjbvd2+SfPYC
xLl3qqnIbsSh+Z40KKVoRAclYu7mUDt5s5Rck31TG9zcWniaGW1nIbwgV1sJqJFz
TMmuyQzPIjmlPjOzBfc1DYFRMMSXzVmnduPPw1ipIGZx95W84A0+FfIGFYRgcNzR
dvjTE4tPvk1LrwRZRIxRHhRYE42B3hAz0zidC1P+TtswINUNu7Rq4/gTJyYACFeT
HeWjYM/x0NZ2QQ8MKRWvEAg1Xy0hhQ7FKN11ziBYm0SngK3X4v53KNQ8Xw/GWqXy
K+P36+9Z2fMITBkguTcKpj1qURwF6R7UHjlxBH8MjuZzKU+vtu0lJHMPLCbvSq4V
r0ZDLIM1Pnp3axIgi8rbBr8R68AhiBxTQsha31KhfLw7ytk8PfIXG99Co05LMsKk
5nDGfz97ahquU4PytU3RTHBf6EBBSn5hGB5w4rQS0I8NQm+4Inlp2kfE3Ql3IMR8
CsHTLmK+hESbdU8g3ofEdjHrBbjQOOqux7xiygPSMp7gZVPhTHlvzOmPPHnn6Ehc
ZuHZiN1hzZyjECNMvPlrzmOe8NMxLV0p+snYNvIVbIF8+Tl+RaVDtGWC1Uqp4Kf1
JOJo1omVhLfkp5QZWIMnTIluHTELRfoPlwbydBacUtyhHVCXbxRxYS/OCkhLZ6kF
43R98S79xc83iACE/ASI08+X/z/yUeZ643+iPvENo68xh1hfc6P9SE8N0rgBkGfF
dfqRAXBxIfsvUjj40ztssPiXcpJIXg1UqwQPMR3Iqz5K32fzN+kr0vEjJlDfsyTQ
sJiBgpIDUcmSEwPINazU3POzqpG6noRrtIcs7wQYxV+i8EfYk1VdkRSF51bByxIJ
9tmFIVwWWMaXNHKCYNBsOwJEJTFmwO2APQ5q0Hnj0wPTN1SKnf5JWNum5opa7Uck
vSfQh6Co7ullWH4u8RMNzhHUlRs5KuSiRPLALTy1H76uKD/Mgu/9mAv5EnkbTz+y
jH8wrig5PPRTV95kbUzWqcHwlnQ3awEaSZ6Tv2a+cWiqCQV0K/B+mZiJkM3x4bZZ
hiQd8xxYC7buYu1KikO9A9v1u882IDu1pe9jwbJRpkq9bcoinob0PDn/PQrrpbKr
k4spZThVkFprglMhW91iI8a+WMynNVv8gUy0/AfMBHKUJRxesZlH4RTvfB9t+Ox3
iAXc9nOJk7cRArZQH/uFpYKyMilM31JxeNdA0YfjpWgnqZnlKL+W44LFaPa2pCfw
F+zQGvuwY+lefHuCUe8itDxm4BL9o6SS6Q6C3GjDnEqmuldG6IZxAQP/1o1yHWC9
7ZnqucebdtEbeqhgb8kTBbSl8V6wQgfJeumZsHRbEoq+czbrufYy+6GxHreis9tq
1HpywcQH2SjyKkgZXDdfWZWfd65EoFvb25fdSZskPV//ar0gNw9+nilu3+J1VTZi
7peY61w7OjosTwJA4NbePpCNHuD/Z4rgvlkeru0gIbva531fAqeL0CghmxDZln5v
RmLFMvUR1bjZCeQxPCG/XfwtYVd3pot8IOHG7TExZbEz+krMb7AoPzVodw1n2NHR
XANnfEwVUTfto9ujTbNak15btHaKllraYb597Dio2nUy2ZMGTuv1xjPK5gHYksOE
fktHwBQHEYVR4/YnRFbBBk/HBU1ONaMFheCscp6mvY/FzdM471RBzkPAuxvUCAzu
f5ZAzmHnJk5tlZX+fsW8jm8iLXvWMf8wUPinudOrs3+Bfl90v+cvy6lMorO3exZx
opf+iVfc+JGdQAKw0/40TTNThyHbF9c7m3DbyHcKquHLSHw5thZU3erCxL+Sgyad
CGhp3eFh5cTBoubId6o5dQgufj863pZmcsv2XiR7y2AaqOhUme7oL9vyMmjsq74V
vgz6aYNVZMrYnZTOypQYfAdIirtLhIiTOXhyUFVwbVMnAA1QxuWHIcNfxjAxvWL4
QXtCkjI5/bqo2eHX7GrRShPp2e77diJKMsHGt0LgJoLWsCVoGovn8QEl7gwN/rxr
QC4qO46UB4LQAqMUDFsoaReifHbZ1iEksi3gjNZo6UY0YuXDT9riZMtYI1q9OPcq
nXnbkNsvOnsCnB8W4NqmYAAEmosHvFV+cU4x7k5FE+hJpImLgH5Oq3Pnp2rn8HzX
wN1f+QlZVy+UocSF8H2/DhN3LY9qS1g1ez3cf3aijPriJcgriGnpM5u3tHCZ4W/+
S0bAobujgH0u9HY90HQ3HovSDIF6TUrWLLLxi8y/i/UXl0lyzNp1nWWPio9z6j05
dJ/gms+Hzmj/LetxvA4kEkMShESw9CZHjslKyOSAWnDxPd2qQRVd+KxNItW/ax/X
2XnApL9nholIkZPa2MHZvLSSei9jGjcJmHdRmBvntUES+zGUCsafONu3plsSaSHl
HaOsrLv/vOqVGmkuuhUwy0vCTGuVcLh0rTidt6HFOFB6+9a0pfTl3TEHrx0y1A7M
1nDaMSXf49mdHe+MGxN0FmqWFW0EQTJSwIlIGgdqF60yY2lj77sfkQc3AYDCDuk0
Vz5ge/coyy1Q9VzcWzE9BdBpmGBaQijS9L8hVpEDEqLNSrUL7vYOaSCzDsSu/wtV
lY5J33IvmFfaibgu4phJ5vDXVgek10Y8sJ/UXrVPk4k3iZzGTNcq0E0iP7MaHpxQ
vbBqwqD0uY6A6IEKBLoV6cxvuTDSB4GOU9MFCOYyv5WyEUj3MsUWR9VbCVuWeEm0
C3SqOYzc39xXi18JIHOsuNAwK5fm3j1QcTauliV4akS2Eozh31QR0mr6TaD3i6iN
wwvwEeb7dmu806OJR5Jn1tSX5WrodTFikBkbqIZk3lJqR9XxwLixzX5RdjvMvV2W
vyujFJQraBZxOaLC5PBT2jj52DIzBe5fjGuPVreKAnkHr95AwyB19mzjQqlVOCfA
2y3Z/9QeDFp0FrLQb3UV0qElJuK2yeYM7u6Skqx1+yj9Ay32fLUwy2V5ChRBugLJ
GQEvXWUAnvrR/+mqNoCCK3IC+axlw+KaanIP5c9Ad9RzFm4kEaD+zJfxkEJrlS4e
WgWqaHylwXqsnD4DY3+iZaWh9dABVwecCAyES2W8/QfRWuNTdF8f0LzkwXWzQbHx
nGuKqc6pvvLFDWW+vUpCetLoRUj56reg3K3XpN+CebEb3P8hB+jduyxCeMvhET0+
0G3OU2j4zoSiq4CLClxMXkvHJEzt2NyKZTZJrrpjsOmje0krOKlHdo6q1axaBVD4
kD318gceHrSFnQmWbqzgBD0ueXO7mCfZTeo1i0FmCFewOBJr8/WsjjmEHF8t+9nm
wWDNz4C9MuRw7VP3RiGjBjgsXa9o9pxarWheyXNq+4EDnA/mLlkgdyNiFwEsi523
eobCIEEQbc8+bRGvicppU2pbKsimL0+NVJhhcYtXTGQadn3o2WdzFWWD/4oBTpt/
q4CpbNSANBtB37Fa7+oMe77s/EVc4iwzdkxG20PiXJ81rSv3zWh43/W653ERoSgE
JI97H+K4ojQEJUkUnujiE6lLE31k/iYId9BoCNyXWmM8xkHa/lUqftoknkbX3Y3Q
PvW/AoqWeeOJGl9zBllpNZqfbp0OZGP6fHCeO0CObzMHY4QKfhMD9S2XFJClO3ww
65N/Gs1Rs17KJ22p5hln3SkrGICiKph3elV145BB89y28VsRfOB0M2HtD1G29T1f
IcaqogM7wFTZ+oOxE1GoE1ie8/+AlTi9LnzGapXiQKa5vKTWyd8GHxmsRpUzMz0Y
Bmr8gfqkGlOtdVfRNDbfkim9Vtv7vvKONcf7LgiwndTbrnxr/uh8C1qCIXcZ+W0p
lVD/WyFUKUVN1NaVnl3N2yYv86H4yxARPvJ6uFj9BMGhAE0ZM3SpUmDDlXym4+Yu
twJqoQ0Ui7VmOt/s7KnpoQuCVN60/Yn8Ukd/eXEtRljx29FVIb1I7MQzOzmlxFCX
b6c0BRulfhxcS8Iev9o2h9J+wyrRHlmZDm5hEDbGEM/g6tvYSoYsM/QiUn8bfKbc
eMXhEJu2lTMU7RwUbaCt0FJ9l8x5FsuBv2nI87gWPHvd0F8xu5yt9tfqmhQxFVAF
NihUhv9Q6GRaLeekoCnM34F3sa+mdOycDU0BpoAcurS/Q8mb+awO/oyWSFauaDjK
004cPV9zcX5SKOl/l3jMG05eISv5qofjO1mKeWeXeory8uKw4qq0CsTNnM5p4b0P
y153pHPga/COj7Di/NVLs42+52NgONX2u/8jEQ0d5HvnJDNRqlGNZmmtoQwu29gx
R/JKHoWokEDSvp8RzTcl03k90Khn/Mx9grxjLpDizuHN33irSpJ8d+IBiP0II+ZE
SqmdWIl3jbEK254EiOqJ7VQrXD4N4WfQEx41P9fgWcHg9VIpyE2OpK6tECpdy5GD
BIF4AI73cV+tgsXEYDAQWh9IYMbHt0p0GiJewuIeaEK/hpWZaXtpQg3jxBbzqJZI
20BIXukPZIvdlM3dz63afRaGvWz+LNqBNB87LTlVqWW2f2eQMIX93LiWiRyyVjNp
XLAEeS4S08IV6PhCQ2qKPDl+JzqYL8Sfi+HtLPAjo6Ux1MPQ3/414ZP9PPP/wChM
CSlJfQ0Qj6Vo1U3fcdDw7VTtliMCf7rO4kndEolPLVccV/BWo/dInGifSKCxcqQb
3zglEVriu7kizR4ZB1KqX7dWm8JMCMr0WmTszpQFn69YI8PHAgG0fJNQSK6a7RoU
j0MUiCymOcTNR+Ase/4wsYY7wUJpvJZSZM9OS6TelpyVWlX4PVt5o3t+UQkmC+Oq
3vq84GIzInWhS00Jny5bWieZ+42W/Tdr0ZTeaDJFzYmT8i27ItGj5QfYj6U/6IX9
+xUjOcsP47b1owmHoWSP/ga0izKIL2w5pBuJ00vtqAXt4Z7rdg5HGSRnzSmIlm30
UcGfnaLftLUI2YHCyyB6N8tAMoufocnmCTuwBNPArAGkRtayv3xRhiRPnoO6+7ak
wGGf6G8Dpi596usYh+JC32Bkw6GTvPQhCPm/yC0mPBcnDCYRgx1VIF568Cxd2tv8
R1iXogkkGP7+tlepEM003NzjkZGXImE9bOALXm6Ssbtvvq3CehMoOzExTGc5B4RS
KnvTcXfitB5O8IoeqZdBgDX7UfO7dw4dmFlhK7fH4IdNcHeiz9kFykppMEa5wcw5
eYMZYAaGGnNo3V6k3ETLMEbiuUBm4AV0Xg6uJFVV2Jib5cF3wEst5oe2e1H6EyHF
OO71ZwOGs1hAGRxChMT8MCC8cp4xZiLpB+NIMfAsTTURv+kkcEDVF3y8oWIZXCX/
tb7XbdjIaiV6NSIPWVBehISHT9BUYu8MCsDK/JESZIUaH3W8zJLa7XPF7NtIwJGQ
ngib0Y0tW8/aPphFS+Df2VXzHvkkMYMUTmyXhCSta+vmaH6CpfcMyKWC3IPRs9tA
rndnLp0Et2Kqew7FZC2kgfWBtvbCci/ve1wqbXIFPhfC3p+ej5VdgE0K9RZII2Z9
WC3xplnxpmd3PlMU57gxD7f6k6L+kBqZp8p+DL3OZiEJfg3Eda/vkvqjhkZmdV6M
GwzkX2lPLOvv00wn0bvw5gQsdEzDmZ76II7i5GjTaFibHQTYKKq7Il2GExnZrZtc
9T0yb/ELe2SMbcN3yBQnKIhiPTOLe+C5tCSJhrTNukWvTTCcu6VIxYaxKT7fW7RM
g41B3P8duVvSRuwMoo8C/KGDiv0/3gHxoZCkc1BqRrDOqRLdHqCpKQHrJKpUkhZY
rPuMeptMGCYjHlCnQaq2JWDgUNJmu+d19XXEVk5Gp149ys79XtbfJtJ8PJWIOvEw
VAZ8TcHSnxWbOWCz+8hNBTAedYbqalBY91rguLWuooeYq2FKVvF1T2A54v3fQqG2
LKsjPybxVMAfLrPYOMKvToBytADS5VqPH95UXUZDpW+AYprX6mSIWYdr3ebkU+DP
rLTtzVOW2Tfkq/zyvcGn5HrRr73tLudIQGPCH3expm+ypkp18xqUONernRaT7LRZ
1DC1Uus5UvXPvlPMTIKsIQkvcxTEsAyyreK0FHLfphw9HZsmLedJoJwQI4PeR96Y
zcWv5kxnOLijZjJsgH1qtwwfMpBzsVu1FoKJSiAd7Gs5JLhMDjlhDoEIADz9hacE
nDCFHT2DWV3yastrQvcSnUZ+YxcmtjoL5yfvtSV/L9Loz8TVShUga0RYOFWeOO/V
NspxxzBFVf9loTrn8zgRbx+eh/si5DyjajPPqhTm7Ks=
//pragma protect end_data_block
//pragma protect digest_block
lARFxky7FMqocKvXfsY0Ps27d5s=
//pragma protect end_digest_block
//pragma protect end_protected
