`ifdef RTL
`define CYCLE_TIME 20.0
    `define PAT 332
`endif
`ifdef GATE
`define CYCLE_TIME 20.0
    `define PAT 4
`endif
`ifdef POST
`define CYCLE_TIME 20.0
    `define PAT 4
`endif

`define MAX_CYCLES 1000000
`include "../00_TESTBED/pseudo_DRAM.v"

module PATTERN #(parameter ID_WIDTH=4, DATA_WIDTH=128, ADDR_WIDTH=32)(
    // CHIP IO 
    clk,    
    rst_n,    
    in_valid,    
    start,
    stop,
    inputtype,
    frame_id,    
    busy,

    // AXI4 IO
    awid_s_inf,
    awaddr_s_inf,
    awsize_s_inf,
    awburst_s_inf,
    awlen_s_inf,
    awvalid_s_inf,
    awready_s_inf,

    wdata_s_inf,
    wlast_s_inf,
    wvalid_s_inf,
    wready_s_inf,

    bid_s_inf,
    bresp_s_inf,
    bvalid_s_inf,
    bready_s_inf,

    arid_s_inf,
    araddr_s_inf,
    arlen_s_inf,
    arsize_s_inf,
    arburst_s_inf,
    arvalid_s_inf,

    arready_s_inf, 
    rid_s_inf,
    rdata_s_inf,
    rresp_s_inf,
    rlast_s_inf,
    rvalid_s_inf,
    rready_s_inf 
);

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
YBY3/CNLmHFvuIO6jh2vHwC8FMjUD8J8Fvb1the6ielDWMJprbAQYo6h37pR6JS2
xS9Xiq0Ctgm/kvFN6CAlj2dnmALqrSwBca8cCi69kSsD+FQmak5dA0FaYqMyP4Tv
mxksPnFb9CNOoOJDmox3CLYiIefJo4aVuBA94Y0sTOk7LPjTOnAwuA==
//pragma protect end_key_block
//pragma protect digest_block
jeha5wX28mGoOILMRrkJW6bf3WI=
//pragma protect end_digest_block
//pragma protect data_block
YgZJfFhjSK9iP9k01iqWyiqkqsyAzUCKcWEmXVbW1D1nD9NLZC8njlaTxP/wEN/7
AL1lXpfnwxI7ZGvmKCzFYUog7IeIfGGnQ3awKoV/2XKa2oRW2vpjl0ILiGC4+6Yg
teP6QUgp7Xrs7gX9Q0Ueodwtl9dL0L/aPrZCO70/sR5AygzIRLH2G/wrbVROID5Q
49yeLiVI51RT1fqZPASl9XPrfTf+GqOsg9D7F87JczKKG52cSk6PXIdB8gAiseD/
ZrCXKwDJ8+RVDRO533tp4jobFfcZBies7FFRpgM0/5DzeYH3COAbQKjRTT0b93N6
4SQTC3Jh7OC/PMm4a+KqNE+S6lfmC/o5Nn5MNWlh/fNx0RExa/RaLp8v3o6IS45N
/VVsoJLw+bH1mQ86QG94oppKwF9Bh1Io+HIcnnvkEh9bgdw4RVh3hJZDbr53hLMA
U1E6I0LuEhKT7Bpaszm22unk9k5ZJBBaE+dMqdtPBfH0jjokAaK61r8qrCccr0Oh
Vfd4gV6blKFHEFEd3PZ0xLyo66sFbJB0OD9jKirEE1mpxW+1g3F23zJ7fF/GxJO9
Aegvd7RSrq7Q2pNWdAkq+92PWWfbtlaunzIGYx6zxgB+wZWeLDJmlwQDjSa2S1mU
2UUMzfbySy6kq1WIxQLgaVRnBbcGbX+hXhIDuTtxyl7tmfJtiNzesi7GzJ8Bg2+1
f+5+/xIgVesEJYXUOby8TfsfEEfzy7nbr5It5JNEiJKaBjNdDhw6HugQAdHZmXRY
Lk/D+D0CxJKhOFVci+g7q6/GQNjGeMklGpTCKAc2+3mwm5MMBQveK0WRMPtqpx1B
n3ujDTJsVrk9PP2hOIUIv9c615CE7BlgNLl5I067QjBG140ieXRV13kFguLE3TAm
q5rlA4rOhm9rPzjmnZc9bOUKp2ek4riIwllaOwVO56wO5LUvt3UuxKdd7Xg7Ys2f
c6XzsJJuLzN+Wo06MzDhApIBZzKTyc9pwbfh9/8X4+2nsO8r2Qb+AY9RU8Wmcr3R
dgb+RFGYnFFndR4MceAIa+4BU0gxFoi4UimdS68R3mk4biSt1pSnQ1v2P3JjaLo5
Szc6+o+9LqFM0m/KYDlADu5Tq+xGdaJXXE66RA54ufDsMPd5myPtEEm+r9kIJJtI
9Ato7Crky84D4JWeoxg9UXe0utKXBwcGgeLhD++DflDgOsnmsYyeSuXa2vgDNfzS
5gZbjJUvgeGRjA4MbnzJ9QG0wJIAbRMHzlecsNWJ07ibOf7KKZq3XmO9lwryNVmc
f9sy1j7407rdRUKLimmoxtZgGnptoJxiYA1OTCQCqBji8k2BQ8vEmqQAsMIHOXvw
7dOk1GsAP/uo9H1XWNV2M46WRuMfFPycMU3gMhtMB4x01No3mTB5UhuSEKSMwM5/
9UtN56TlKjFLpcghQlv4JnXmVZI4mx2XbCp3m2D6zKEOY8fWfLTmIH9w3C8huLwu
RrGSSYvVurhqyU8e2msWiPARKA9BrRv8g4TnSeZ6rJ1AcQc5yJahAUeB0Hrc3VJ4
goguVsFR3Y6HJ9Ev0jnqx/yUvd2Y1315VaBgz3jYsE4TdUOhTEUbihjusvo153fd
gFj3tLbSQaLI767BnAbgDsN8RRzsJfUHE6JOs83bWT41iQfgdiNq7EhMxsllI0rD
ultx6akAXHDaNEReSSBsG5qeo/uuA/c2YTVKmQoQO3gcAJc+cqDAL9nmFZai+mEJ
RfFVTGTff6i/BSWtsiR4V3nCr1rD/xvalBxMl9/dvWvgSzUZFRy8IjYWxYIFt5qN
7c2RMEdJ7QRD7N4Lekf7ypWS9ApBYglrd3DkE414/HGKWeNLn1+wopJS2rmnAVSH
BB0YElFIqt0s8LBkSttzyvFA4HuNRe696UmN1LcYm5FHZJtCcT/jLaqXZjhIB7gO
EN7Z5olN6vIGFpEEdWEplpPQ5FuQpupm8ngA4QrCLMETjG8wtbWF/QyaNUnfjjmI
Nqe9s37i7gNeaDLExEdjjicCbmV2DRX8xob/zMIrydTbE8HTS/oGye7pwMVh3GvS
pzV2+GkYh+rk0UCj+1eHjclepwPC41tWKIxGhnCCmJ+HwIwkrqMIiNuVGIYcw32u
N9YJWsaVPSnemF6vCiHSZtSCCt1wwf1DeZCC/PnycRso1Tyo4jsF8UqgdXQzv7tD
c8Gi4ojARe6Bs4w3vrwiYd1M3Wu4Cs9MMDZF5d0VbvLCqg++6ZVC5PjgP31m3UOP
NB9ZpNfIQgrpySigjf1WyAynIDekcMQ+bMjf+ctN7F9J3j6mkqhdgquXnvi4IsQC
ZDq0dgNaHTfT0xaOWzX9eFVF3U965t13UnTqYx3LWd+ZDxgcz6I1161tuPu0fINe
RSv45b+AwtEzdKG3tpRJaH0K9ONzkNQCVnRfAK+Ekm+ffCmc0WbcMXsrRr4BmPx5
ctGscJY//IvL44yPkmajHmRTUUlDtG5cv1t5GzFLCRL2mz7NeyrwlUOHgs7830Aj
yCL6X/gXqq7WC753K6tpTUSsXtJjUYQ0Ho5RHtL5/GvWIx+xkvI7JgfNmXJNu8VU
6B1GLDPwC6OZ6gQGZMGCCYvYCpB+vV+4Yq3dEByqkBfBYAcA/X9/Sie/9s/EnKbm
lrtGo6C2km8v3R/NWXsYz8x5V3RNst6ojZ2gV+ekWEBPOmhZpTGLnt06UhVHKdR3
E5v9hORAvCVUonVTclDJDZ9HHLsaZeHXwIgLcbi8LGp5o5oW8QnhdHI9JgR8VAC5
6rSCdja32bXu056cTP8Dz69Px/67Oj04+XMQweyqDRdVZccgv4wwgNdD85t/m0QL
/miZ4hJoEQa6tl57cqdDWmHB56JmSzgQ7EyPw/n3QF1iVl9mpxEuT+lq541NSP2+
X8TIvU3ZWUsVvqf10h5e/fs6Ajqqp/+hdFGEC+PhICOM0+WJgwhkOMUTIUG//OHq
aBuYHxfYKWJhaJbapMxOO9lL2cFsVBaSktZ9CooHluWMANwjCqBgeUdL76aYI8u5
ufW48K9TCIEQMHNVwzsQs2E5U2Jy0L2YKfRZ3Gkuv7zaGA6QHYxcevAxdGcVo0SO
TUVsCPD4mtcJdiBHI9VEnaIwbThj5vT7PKzdGUI6iuItzEuzJUc1AFu44LBUQSPi
yIwCEv1t+ucHjH7dFecs+YyUyB49FTS/VjXnwyJpz0PoJmLT8pWGa6GOxKEwKmyP
830ZdqJodQl8v8P8zc4+Zr7IPlohGfX4D497FhpFWoBzqeRewbZYngbaWjByDTiR
9X4RZIgBLfvVcfGlSLdfzkEx7FtP6haaZD9RGzWrM66f5Z3JW5vS4b0FxV71H/O0
GiH01XRys0FW2+A1DDqftz8oo4EADXZW1HQVp0w+aZyDcNbkhXQubb+W5nqqUubv
Qj30rAtH0QAk7z0WPmXWDAANZ7Z4vyS/xSqnAKBuN94+vmVagomNfrVFSYJa5lui
Shi0zg93FWO5i6VGz8TnkXQwIAo5AQV9ROCNXqphC79Hr7C22DI3U1dTkvyxCmCp
R005/T6hDumeDXGTpDX8LeD/YLMBY2j1DvYQ4yZEva5vENEtq2R1q7aJEMW5UvvT
KdpLmM2cMAU00yv2PV1powU70w9SqW9S7AqRrU6iAtu2wbhMiElpKT09YU2IEiej
waCk1lI86tDTTxpBT3WosuSe1JuIBBlk3/WWcLOmZiFaogHpNtR/MTDEtZBaXNkI
LTRIKgr4Rxyakecocpxi//uSTZzwK/ImFUOttQNPkGuGMFND+w/sr7TImc6ewCLe
U24iPm7QytVD9KgEQV7GtzJfQVKS0CTgrS9uOKz7pjC02SiPC6ZGOs2JPTNQUga+
ibyl296CPHp6BIFS/uaYtYJCHeYyBWn/dH32kZh1feWYSD8ZQU0sM8yWcDnJdDNQ
VF0h9EG4nuv15l7ofgI5kP6sIphg4mZJo6agzufZpzDJEwqjG9H30rdxWuUZzVA2
n4mkmpVjSUSrpkUjn6zKXr3LZyqpotyXhytrJNGqxtiE/Ae08hZ7i3gbC1Zf9mfI
LyyKnue8y8Mb8eUKJI/1zl4oqTfVzBEPL0Qyv/SRmkG8Sy82ndGY9706413SlB59
XkTODMtV5Sx94EJQ1enri555tajcFLKLwawg+U9dwqUEwrk7zLI+3JmhsLH7Z+8O
AFJmQkKnmZj+0Dsp1nx2DjrQLVBIaqLWljjhaZqYAybzLABvc1qA8Zolx5F5Ej3Q
vTxa+rjAXHbCyLwh2uXeZuE0tDnCSrHxwFrS1Whwmo7jVJlCTSKuQXRLZbsDIWwF
6RaSsJtqDaaBaQ8eIweHib9pvp0TShODOEEPBiXP/c9t+FB4YXDPJMictJHU1wGs
7y7T2ciseJcumWYE2XJUmM9ARGG6gwnpbGz91jHAet+zEc7YXzVUhtzD/1saT8Jl
yYUyDw9809rO1MBvpRC1q1m2f/IHCjBXIIk3iwglvR7AbkY4q611IHjVPVoXAjPo
9sHy9M6jFfO01t5J7xoacPQal+0m0raEqjYvDWziZ2TsFMmmkxN+VEYCGAO08/TQ
C5z2Y3v/K1BmuP2CBYhWf+S7hzOfFfTRDOOoyxQYthTZP8Jo4yGdrO9HckqH0u3l
+J3VZSoQYVao5Z+LZBi5sHW/qj9oiyUnGo8AKOxAwDqeAddozPruQOhdomwAni6i
anxWoe0hRui5tzS4Z4o7GPNMfmQmBrOfNcQx8F6c6BuHosGW5y5796baDFBR57OA
K/8cLgmANhOTzk9JrcXy3A1TkbY6nqv5npPbu41WUsdzCy+VPBNRR1dhG7u2Pccn
MVKYS+k/kkBZQcwcMs5Om0UAavXO3JIFn0Nx/SZSG3tYzn3cMGKLeAlmWpS4w0S2
c2VnBrFCtaIP19eIwhTmU1Am2G52piKLMnjg1+3BNRumqDfBRxG/3QT+YbbHvE5A
uOxwuMHRUjJIQnVgTdBUAr82+ZaBUHZAqbx/FpttTYGeL56gpz095TLrj/RmpN5S
qU/ZbyuXxM38AkuySnxPT+pmP5MtVsXowRFdpNUSgnq48vfYaTCTdtHQXmnAdptf
JDxNEfMQUp1UAjG3T9T5USQLvS7sz0VgbiZlFEkPZtI4ZsFPRFlzmu07VN0zuJGK
SOiIkihMtqzcu3aBR1i6EDLIWatfy7W57JUjADYApWfk7xuEXimsRPq6E2nfQV0q
z+Ri31HgfUMaBVO9GhLT85lAxSVNS+fRwigIPIrxXE8Q7FtOVPVNrQqUiYPUr2k4
R7IaTalLVXc0WgrfuV96MkJLfjQpdfTRrcIzlgkbj0xKTJukS9t+RflbELVeLaAM
ZJG040t6Iu1w2nDYW6f2Doy6qxN9CU0wKIyyQ/W74a+3JNE1tMn2WsySkaif/4MI
y+W0TMmDX40jcSn9zgkrNG33Z8XLrrGijPx9mnyG92dOG0G1MbbBxkARvWUMkMpE
gvGPD+qf8PIOCDcX0bvIGoNqyEANUgz32PFp5GfBMFyF0RdR4ULp1I1hUERmuReG
58eWUv2joDX9H4/884LkEG0MclVekl7I+TjlDDXK66O57WQzDGKpKmcWBDLAIbK4
97JSLCcbwPr0Wxg+/jkMGVLayLNvZ81NgINC9qSXQDq2JcWzgh9hZbRzI/QNvknd
RswLq2swIut6P/SKnk1rUCps3EI5lobKGtaT7U4pqFHUwrXp4/uCruF042XQUFfW
vnu7qy4mMxkqR9iOs2M5Oz7kKRrCmeHqudrZ/0oSVXvbLUuVNAT3aZavudmtMUCi
vTkm+KAbdFXu5SJEE80VBAnIXVjIuvJN5IlvUtNvzjCmT1PzSv5kiBfgLgwrtWdQ
QFopgNxzWq0uEzTFbqp1pp3poqM8YJ5Qh+QIGk1pwYuuJ9Opfysm5CPrzpd2pxTK
CsARxe5kGqjiy3y73pvfvJKhcHFIVir2OV+jcS5At9/bnT8fOzz8Za6Wkw3kRQpD
ychKH0adXr/YsNsJhQaSDRf52Pt2ukuHqCUcid57L0hbX/mcu3oGR3EOdGngaHVq
GCTO22N7DEG9gTT0MqnoXT2m/XXIDvNgyObipyTnNHQrsyiVg2zj5Tikb48+Yusm
zDo+uvlNOAx4tHrWFiEfJToa4iPUGV7mnOxzhjyOZDJtHgAuRr8JJj4AkU0Q9Kt/
GKl/lBwCyZLy1y4uQv45wrEQ2N+gWJ9jHuslYPuzHCVMjMcIsGrMM8aeqKi79Ll7
xZ5x3CCQj1Pw+B5mheV4xk7z8xrNGdHnIFgc75tLaFgqMLiDSL/Yuclhk89wFLHF
MNfbA/gW1gOqQv9weglb7CMpBX1yOLtZ9+qW3MAh75Nb3PKQ2H8Ei8cWJsYY2b+4
sR8mY05UwULC9d/qFTEUlUAM3yeHhCTOesb3GH4coXn8whAXmydH5c4BneftQdlq
+lJ9mUG370bqRwRQFhABb3RG3H9lHe8pAfmgDUsLG4V98ZlesVx2w8gDWw2/l+M2
XvkUZ6aEYJBIIJKBHf3mzSnhHvQoUps8hXytqfSw6/jFufYzjpu2XMoqc1HhOzYT
sHWB6HFfOJyPbV8wwYNqLy7cH3GjYr+Fk9XJTjiD9lxS4zloqU0ZnB2cMSWtvl8L
HIBQp9YucrPn785CgTUZXiNsnc448rVKlwy2Il8qKtzpU2e2a1yWHcVcKGmF6HFZ
y8P1WvN2VjogMFqXyObXQsdpsp9LmZ9QOoP4XcG7w6jhjUCUdHXufyUl9JnlBsC6
rkC4vh7CXuWQ8uh8AAXZKjPZQVRtnBBhYXfFIOqz4Uuft/2z6wsY48p3Wj6kxD/o
pdF/sgPMQy2mtSIVuHNJ2lYalU3NcL/oxEANXn9u/XbZmEQFhkeG90zsc4yS8l0C
YbD//9GtGWu9NOTNsNB7z+bo833AuOTaMUf4Vzjj97HwL4swp74dBEnMDmrqxBu4
EfHgE5rExAaqrxcd012eUtlnuwsAshwlY34wvCVqS0V5igNrehK04M0Z7LJnliG5
+smTieaytQDom65gFtsAefv8WZ1yINrGKOxu682BcgQ3n5cIl33gt/6zSeDR90JT
RfaMBE+yKGzZ/vx7yuZGzcjJUPGqA2nb/Lpkxz5L4EXEyd5lfpYBQcUP/b/78oYw
9EOVWj3vPjUwDZelshik23JlJXjrMQUzAe8Q5YWYdduILDqDMNwxd8E1V+R9X50F
qT5XuUUmm32m0WYCoGCyg4rYAjb7U00Ar5UOlPjNk9IyaYTNfZLVAKDM8D11WZCi
jPto1nO4Yn6Os+ks5DxCglmncCgnFNO7xhFhJj7tEEqUdiBVrHdDfMsj5altxwKQ
z9OOHJEHF/+upkDADeGBTPe276DHYttPBtJUremxkSVzqBuh0WWwyS/Ng1oN9HRF
QhRGcr+UyrGPNnvLahWojRUsffsDx7JOgY0gOCU/fHie0/TPHo4RAf02BskwAvGB
azDzHAFqFUMtTSJSo6OBtZvv1dnWnwp9qFUmmuQsBp+8iC9Fw/k7/lAy0QAAzya+
g6Szf8mJUqrp+Tv76VXq+9UIgnv3ilRrDqPFLE+iPbffbkBeySEJ6X/cNKGFx5xe
oPUBQPqVE3GNHm6v+hXwJLkhZ/qq3M5y128IWqDv9ip6deUot112NOGQDP+XZpvl
qfwDza+trBdrDoBo954hhRbxlbdodBKUQybSitPH0eDAE5xcRu/FupBV7x9Ye4C0
taEdJavbygGGqMb5XSxSUSMMs1zdVwG/s9/SL64Is5RCwQJCqEnAyN1RboYp68rg
qFylULJskHEVIvRJ14IPtQYUHSkTUn7Z2Te1C2bAN0M9nfnEwicv9YorQXAzMfQu
0n2PiM1Gumt16W7E7nmrCo1gCUHSPqWCqex20yfVh7rFbrXrDf9SLqUGrhdbtpwH
1zSmlzsVWBRj3rjYJwEgTGeQSK+cFqkRdvVSSd1BQQTGgtb7PznjHliQzdgLcQDa
dopTPBA0Kkei7ySQFbLWLbXEOpY/8SPQn12RwXpm6fqXMAA9Vq4VgZKf/drP/oAV
shN4q/yO60X71ETRtUIA4btx21hLdEFtEu1Dms6LdkM+x7Y1dTYzlqu8ih5Yr89P
CFLywRHDcHWTwbTcE+COjkg7Vq9y/aq7k5ZRU1+PP8TLH4+CbZg2SNbEWjnmJr+X
ttPRZ5dYceXcZgEkZZZoTEMR5KGR+8P/o4bbX5jHHuXnq/yfkMQ0OvSjiz6/97a7
3nIO7Q/nvs/jC29BpZPBTfrlLqaGAucPZ0d6ceic8VWZtQkcFmDiNI4uVE7QNG8S
/OceCS+yEqALXqsGppsAu7aeits/+Rp93SOeuhHGGYushmVb4lNM4eqRNh6il4ae
0GExPty/PgZ+tXN0PftV0/teVdjleDbhFQZyAas97zqlS3N0nbRAyQIXjNeXOyas
N/GNpHgYpwjgT6Y763dIXBJdZ+3cvFTB1CivhMAFHIeZINfSb+lxdagIv99eGFyC
ZJqKl1Ya5E5xEVWS0Mv660ZwMXxKLSfdQZR6UQ4EO73Fjp2nv5+k/EqXwX2at6W2
xuJEPqINtzVsBk6Ypd1xqyzH8xLFKPb5prSEbq3THqI8x/Fcyo19rzQQWNtII5IB
quUnG2FlDEy5EiSkvnHiRfT3gJV+YloZCKbrgnCr+fII//wOcR9488d6FKunCErN
XEBBc5XO2tJSdOAFFuX5lez4W/VkQnrBE4OhgbffnVxgixmNEY9HLcAb/KF4jP5S
DZZmb/uPBta+TMN/ex7fyoBM7BQjo8JIe+iPHVz2vUCQ0oDRs4+fQk2/EUUDtsri
VQqMX79j+3T2WDkgc9IHsVqmW8PUIh8Ba2T9BsTtVy0SqK410BhnBf+dTgnCkDjU
Nb9P6A2Mr4J+NnX11KZBstELjUck+tBsL7w0R+1el9SKIGQdwPC2uT5lmEqM3yXx
5ctwkaOuzdHz5TQLeJ8O3mf8NzlITrOM/NTmFKhjEHbFSlQ4xGMGUM1A/5qJv5Mp
8WPTSbLZbm+ueE8nv/LGr+Msg4yBSwndxlqigAlS+8CTjSXgNBV6O0OVRUq/yQoF
6Yd2mQuitQLdBU33V3HNGvjSgykHO4shegDVdwXFIUanE96YQ4e3vjby9bIvKH/8
x0UEM6xeuKH2ffXXISfc8WWImlt9aCIFudb723S/5jL/z6eA9mO6q5ietK+QNkNs
eV44U5Tcup+zuz6wLQvB7sTT6Suu20fSXSVhq+ombRDzs2+lJ+1QLdrVXv4E0KER
8xqigD7qkC3qsiBp+eDR4yW1U6cj9h9A+AqL1W11H8nC0Sg/6vt+C75YYAvJ+nZF
nzSq+XXiKrTnSQuw4A+gx7JaOQRC49uroALX5uSQutZKk/UmUWomIF1nqifJ1Vut
i5q/OVGskfdvSSFFjDAdRTpAcfgqMTaFRooK94o+Gy+eZ8YDLAwoNEQIjzWZ1NJ9
mxYz5XjX/YfyL2bvqH2XNikUIDGcHCYaLEOIP2gzwxYGt8SKeZN/pUkNj92p1ctM
HcdxvVI/sIDJZiAUDkamXozJqOGcMe87TeUuZPADLAMLuPOvUeO4pGIGBNFRgHn7
Sf7j1ixprYVeFyoT8jlKhQc9+Dvopc8yRZffrcS5I6FNfBDvcvKOTlUT9URp38LX
BORsXy2uXjQngFMQIG8B+b/6THVdjc4aPDN5gNKEzBN/g67a0UNKW7thfXb+hllH
Tw86yyWSy9DY2IWmBEQ8Tvq5m82K3fVvLOzLSyZmXeX1IEFDTwrIGsJgeJr2FTHb
US9ZJMa6oOTkNHbcuceEp6Ym1fdXoWeVxrRIH1PLN3vi7Z4xYFASefG9gBxzscjn
9S/3qd8aGMGye93nXlHYlxyaQEdBfAvkRSDkUccXg7km4xncROvOvYAz4RqUdDAX
wLrd/OagN8NRzLlMh6IFI/pDJSMECUJJCwJpSGvI+L7j+g7owLtkm9z6B9IxHkjT
P039ph3nYAn1v0MLgIflBw4dHw9MPM+Jbut3vA/dOORD5iPS3FLqkfHS9iH4H/Mo
7C6I7WdnK94dayi+tnxW4SMK0FIap1C1umqWYaUV48wQY9GfxzdQhEe2UzPz0hAn
RN4jKABW1peKdps+ToFS5q7N1ItK+jytfjKNHf5VV/lpCgZvMXO0PX3LGoErl1vl
OyIBTTfOgSlj4RGNZX8g5BWJxm1SmQz52qSubQCuI7VGMNwIjWZUgzffgJube++J
VordHfJO3KoCzyJHhvROcrqcIkqoRIwCUYAL23gEk6nPJSpuKMajU8vZR5r+l0VA
VY66qp4OT6WYbsNhKLWjCDtfkhh09ndvXIs4mz8XoMC8OJo9A19PK1GJCN3X94A6
wffn3GymYo2M8liDPgFGMV0whVONi1z00TUIXMAediSj218u9rwBETe7r0xIRVVJ
a/ZQFGJc741UjLdlL8w1i0jdnNjKO3mpSRvOwsv0O24nDMq/ok8y6PHp90SjAX6A
qq0yYAT1OejDSp3PWSgaRSxfmHeyIhbJcMiL6PrWw1e9xz9B/b+o0s5f2GWZNfYZ
aKT04tHM59FRKOlVOq9QOu2iEQhvYqRjeWkylzQYZF8HzIZvyGQGXJ7y0Wo1wTX/
/wzH7cIaMHrzshMEPyyYRyHN+Fpjdz3tetqxoECOQ8VKyShWJSb4Al2kZOBfPGA5
J5mv6VrPWSBu4IIw1dEWwsvGUu6UKwuPL4P5eUUDuVUiPxSFR/32OjZ0/i5kTY7k
twfNoCAVSMob4eW4wYBviwOLdmUSR23PW4t14RYh0mc42NxQIWR5nnx18eF6kSMi
y/mOzwUWWyiP0mlr0LdYPZi4Vv825KJK2wOcENkja/kyei5++6IiNZB3RySubId2
VMUUTHVVXibySygFbhc8t0gBAa8XY+0s5xL30QImunyljdDwW6wOoeqfRIhlMMP/
3cyKSC8V0EtAiaP6JETRXZTMsCxORC3Ej4pAtxN8MyvWf24D5713ESwXfSVWI7V1
hHfDMOH3BnFlxEW/OfSCc+kjuZGWX1Zy3T2vO4Xft2lvxbBNl7Zd5lRq1/fOIHq9
vYzFNu11FJhAqq5FhIZ9U87pA9kpXg7b/aUEpQ3nD1nbGSfQkB+u8c0AkM5KQWlL
4yoN9iTXDmUiGcJ/KPnqnOjXI5K/ss5BtmQi+Aq95pv2tawGLv26rrx3z13hpFYB
yKfUrUD6mrqK9uG/4Qrdcswiqs0RbMuvk/JfDO4FbHlXXuVRU5mjYGn0NQnRvTsL
mqTX3nT9SNPvuN2IkxEiL4J1ybxfK2VY23VafcGPDKpqYX79ITsKNZLbwPITwhOu
X6ZGQ87Umzf31qYVlYQLEZNMxxacf4SFLTU1Kw8ASz5M2JVREEpwMpRmGgwoWzvT
BpIGAzgfkIdKq1y59Jb3K6536uTvQb6kPsKgmVgASNVvIArwRNWkBUszagFSpzdL
5sCUXQI+jyMghqFAd2VVn1qy4VwwNx16Jp82RI+cnRTI2ZfqHrBBCJ49Y0kxnb2b
mfh4f5+OTkFE0wQYKe0GG3RG4RcgeA2O780r7g3uiNuQekPnM+z8kkInpydTBwZ7
1UWOcNNFCQB8hywfIUMo//7MsPA4wsdwmPpMxJlGhA6S3fSSUaI3rJTRNG9re3lL
Y4EQV8PGxewsQKy1ieoUQjdwNVmNoAxwVyZmQUyp3dCvw7fdj892OVErEd3ZLQzM
Qq/YjnvpaF+DnYcK7hHA9WuMhvkHH6wt/v+80ZMHup5ILamrrl+taNxBVLiK44zO
JdRbyRDM+fJhzi5K/84FGnpdALk43SVAs42KC/b4qCV+b+TliDSZdUXCDS6ImcqJ
rFscjumO4PGUC9WsUP4spE5qA2SPf2mkewAVg4BltETzzvmNKk906vp7U6Ebqon/
6fEAvlccUNKZ2eWoDfzwjhPt2KP5Pa+SihwFRBwhAIZ0K33MQDuTS3cq+tNxcLs9
pXgJhFUCUdyvKuRBO5Ogee8UuEkM5l2QvlTAwXxt6GBGE6V2Re/qWnU/sPSedOvV
iboI4oWTzQvs51noHh3kT8dc4fhi9p1JfZHmsHaf55W4+OTmK2XMu6rVvn1CNPIo
nNDiq8iB8dMcqyGprmk+iR8IMVMNkMrkoRC9SVCnXKDWITs0bwYySD/f+LqZzmpv
IKTK43hPpz1jg7QaOWu0Em/Yzu1jii5oRDaLLHxwIIGZu3z1Mkfn8jUwSRvy6dQa
xV0ezT2aAW3zZXBnZUrrt/pRe33Ii47bWa8C5g69MgIESZZN5ltICGLgneBeOQsC
bnQfukQwfAi66AMIW09fkxKsETlNWS8PrJJ/TjutD1sN8lv5SIz+3mBaKsBuoVr+
ouLji8uBuGks17xnXXp7/mcAxwPUOa75y4lNcR4lqUzumZ+MnwTx0kECzL9iliWI
ehYe9E//rXuA3GyXvKYe/+a4jcypB5ba6j5OZQhA5r2BujjN0qdYglYnDWFYPqYs
0O6xzqdpdZkWfvzPBT4oyVc3xNTvJZx1MYT5na+ztWFFP9vSTFpbuNOGUBrhI+xt
XqOJN44H7D30QRFjE0wZpCiAMo572bVG4VKIhmy6PKqEQfKLytKe0AeLstCQrRc8
/0JiWLeyC2xQQnwZz2voVAkIfQSpYvyK5HY2mJ6THESFkHo0JeQjpdkeHN5ti+ex
PUt8ICMdxICzvwNvArUDk2q7y6tc+zsHgBa/OH6Nwwofty5ut2ycE5KdFhPl/gHF
liTd/TGqi/BzxZLPpL5Q1jmHKmsawjG9Ac6Jy+zppNS19M3Hd443QX0nFQOdywas
GyI0+hl7vVwpgvw3WMJCRW8eUhpdMXmsU4UsEgxBV2nGeWQkruad9htiaCc/DWSz
Y0r1TNZzjmKcOe8GQ76lrh8qpma9lIR9kxHAWVEC4BJ+B8U8ec0B4dM8UpquPaRR
aWz9hDNukLhmCatMkx+QGA3HXIjOjoWxQ82nBHQgrouaAgr+VvJwrozludTiWURF
eDxg3Hhc6+DHtsu1CN5mGdTMcIItl/Akp7pbZ05Fv3pyouLVBs0Iak9HE4O+EL+D
imppN1GP/WeJrEIZmqX32hEfYtOP5r+oLaQpXRjaLbumY2GcNobvUgx2LvpgNTFD
U/y7gc7kIXcE95AUUWEo1168SsDEr34F7My4LPN2Wglqml5V9vnfjmaCZeqjDoYv
L0kvZQxI8m6WsNWnoYYmSdXeSwdNqH7WOuycTVPVuN/EFegP4L8EOXlorXB0TKw5
swfuEyA0tzTLsbzDcRY45cQS5AFVgz/elp0EmMnRZScSgWG0EvSJ0XNQcT8ptr37
43Q2g+jOcPWjdON5u8aEoKnrR0Et+SjWJ+lbVyxTgD+AEV/4t038nJ2BLULb7fza
rEjlbHOZYB6rQZvsWnfbsaLO6LOYLBTegiFy469jr/y5QmYB5mow5jtHMCUPTLIY
KnWrF7zdH0RXFqHpH6ZuqknCaa6R+WcxRZ7ewFNHrZJnKEDs+6ZzWELMOVRkUwKs
o9pE4Km2rKH6WBMefHdPeN1TG0BPefy/yPMCZqDp0zVIjwvr4ao62zkKIFPcg8/a
ud09qTZFzICS0zJe/NYx/JNIfnBAPy5DzWLHLO9WKaCU2iCwcP4Dy2U4SZtIL7T7
WcXYUeYizk6UL/IY3F8Px4yXae7pVcxlzT1Vo7jK0WKKOvxPy9Fd0wK6W7JbKK87
U8stivftNsQNBV28iKlHXb/prjSrrNEKCoPtqQjkn23G2XlCK0b2ZBE8ZSAKe3KL
+uJ5o7EYcIvjDGTbHCvPSGGv3rR9nsrXBbc5qSWzUqPIUaUTAVQixTVXcLvlbQF7
i0SuAbC+OcmBMEFdQa6yYKFNF4XLB+fP40U/N9XhzjUOLGrPK431I4siSQmV4x23
c5xNjWiMf2JtQIDQfg0eWStHhPXxdFZE9Ti0osGwYYoyvHNnIkSgR5xGw7y18iuY
q2nvzFHjiUvK6Cu8SKS2ZRsnfHbBfLib5Qhr0r8YM5brvQa+jfH8PdDzWFh9w18w
rBdYlAjlWRWRqyiwylqfsQOm02Ep0v6kGxDsvK00xvbAnbY/ZWa4ynyFEEz8hUoo
8Pk+FOSMvxG0C77cUqS6mivUR14T3qiMfldW+1vCNFMuWd55K1/aZ1SFiDFtZNwM
wUIiGJOrWaDyyFmLOgVo7GsXM7nRXNU9wZgIZTxvmdr5Il4G7I0ZUSccrHTqteF0
rkuiH68tu6vJMB7UaBifEhh0E/aks5oFmZWxYNODPU2HNpRYiEDsdcSxMVrjSTSk
GKmjohVUT1Xc1PUi0u6xvZKK/1XUdFvp6bHvQd1DzBsgvbhxsW7+b3GtWamH+lEG
bDuPCJ3bqpO2XI+uxZCQONgG6G7qsKXfWDKw7wLne34tVeWtN5dZSnIaYpiTgp6c
kxiDpxrM3pLe6fFRJOD1kR0CM6Aqpl3stms12g+Ix6kZaceOXCbZKihsP0Ll6+yd
GTCmFIFJuGLQw4iWXyzT5Wqyq3IGA1HUQ6s+E5B5C1BNcvVh7EXMgKgk1RB5Q8IL
EzOSwM0xPEl7pm2sBusKBeRBHazY6jYMlbDfTTBkMGcrk61k+WEsOISzLPSOp4MC
Aaa0KReU0ACN3R9zhHCPJuzhbwjY5tUJ8BC8+6FZlL3TXflAsq2fKdaRqpkMbswA
NVcFvLPcLUi1USlCcpBa1riiNcm0NH871sJI9Mgp++dKV9gI4Iz6H9JeZ22jn8Ph
kubbrPjz1E/OTkRAgzBHkDsbucoT/VeugiLhMb498vRvcqGCKe6rQPRo5JaylhCC
wA4JTunIxnPkjS5eArYUScXhIV5w8FqRid7tleQ5ImkMx7fxBNsXIj79miFRTcg/
CuLY8C3oS2qJjtHVkys8kxxv5WAJ4p+qNb1y4d4o0W4SHCpUqeH/HvApRJAF3wkw
Rh0majI+D1+wFy1piesoR9jg+eeolR7G3GvU1bqQQqOUXkOyz4p2qj4Hw99OdHiV
pTNc8rsfgj/VHuB2791Rm6JaioyXwMGRAWRKerSDW0nTMtI6S2ZjRHEfs+JQoQCC
03gqyTTbkLpfKIVFhdQzxVy8EBlVwUHXFlGSsOzPmoWxsIq/HqRvbgn+Zd4dRKrf
4hR7tc1wez4yzdjpSWz1sDz10q6nB7Rkvqm4Ulqh/SDb6qjPhurHxZGvXwNdQpBS
5VEznrIPR8SsvzYfpXnwy5DOm5M/Lwx8pZzF6OOLU7VlwK01vN8ygSYpiCcxYhly
v0MbnW4GZKPGRqB/8lgJdZDRwZ3v8uhPh7j4k7NdcLvU9HSSCs55P76fEFd4n3sT
jHbET1GLuhZepXpyhenHTxBWKnST7XtZngY3iG8peYZbxlm5GHPvzKiZIV3zx64a
edHkG7N5S7nHLyDHugK877f2UeXV+E0sdkbh0eLGzXxuCgzCQZJlMDAJdaRL9yAM
lrv/pqvVdG3B2G6X58IA8o91Xx4Lv4ZOkZWUOxxzi/9C9bQtToB/zpGEiyI6UtEw
F4ff73jqyJlsaCLuiG6jqlfEcrZqPdu3XRr82oPTmJGuVuBKL9viUuk7d1idW9c5
E0gnKZO6ALvQis4FaJm0utIEDnsfDOSpTom5pTtUuqBjWfV6KpvL6pHqRtlLuDl2
QlbZjdTUP3HX16ptGEBYSkkd/1cc8Bg9r1AhzYUWYh8rrN5yht9qGCGNC98XsFd5
IF2YxfLS25U2rJi3+gKOdIyzHloPx33kf8+DtwurHiOXH/G2jvMNQ4B9V4MW6ser
eJ69pu0YMpJfmyJ3nSTHSj+94tGQK0aEjiUO5BUI+mqUuQ7Rq4ptEhl2EsxPrdoL
2SIV6TULb3jQUc0yKd3hUZFKSnNiVYdiTD/Z/IwXvcK3Cnlb+cldkLOmiQz2Rri9
SS1kZ7TuKxcZbYD+7H2Pki8BpPz/jpTE8U2LOzoLbPaDmnrM2FzD4+47mh+qZPfW
bTLnEgdM1ERIKbGZMDzsh4x7camQzF7DmYHbMSHGs948kCVzsMrQI/zS//DdPb5d
q6C78pDj49H8fBdr9HiywQeW1u2wG4nYEJ3akb24y5KQ4NkUQjeFtcCjVozqgDiI
bbL3HMnQ5ymA147klyluvQPEHFe6Z8oPxHIH59aWx4WeU8/8vBfBfBnXOE0kpsc4
CInRjQ6ju25JnjkozKNH0dohHfGLZie7zVSwY8LZG7Y72oN4IpHeC7iqrJNesexi
ihn9NIDPVnkDA03KkCkDwzAvm3tUXTbjF2tTKj/RMLBfkuovpLQBnT/lQCBpdyNd
wEb5xVaCw2SvbG9DrUDn5vk5pq302xbblLwqS7HwlNjMcaOplXJdrTUv3GqpCQIg
FQG0xgqn/S/y7pETj+c/e4fhbrJhvR3rD96Md74uVlFeRrLmkoF6fsdFRm9Iz8nl
6A+i59lm0p++GgfQ944beuZ93FFA5uXC+NKbHrErGA72/1dhfKtD+nYwSu0vFUY+
SWHhtmvjgSIqluYfegsjqaUoYeLZDaDD/C9LYl6ssZhvUgm3aD+yYf4/3qkXPZXw
SmXBxQ22f2omFNP4Sg3m1+6twX1bLDgX5WW7ZN1RQkTZ0big9p5S9Lku1sJZJisp
KdbDY1ZngBaK0DfQYsoo7UT6CsLdGCAKQIZEhSPdxGipJiGJx/n++8mGI8c9ydeZ
FCseNxNhHDY6+6EmM1Qx1yM0F4RxP56+DXLxAzx4l4fC6SVjDsDRDuRUW+xGz2tp
QD/vPMl2T+1z82jU5YjFk9KAG5U02TYGfsJd8WI5skmWaSHx2pvWiYymH5kIFt6O
MuETCdKmra2IcRcvH+qN7BAr9WWprs+T4LqeBjk0u6KVNlrBhYRayt3PGRETDFDN
QTWM/AS5el4MJ43CiNBrGcfv17k2Wdy3Ojp0kthmaM9D42R4Z2KyeVEzcHGPpyRW
r/iEhOsNJMc0EiRv7RtKRFCHB+5KdXXlFe12G/FjLmKZTxhgB1xHdAK47dE1q8ip
TC3wdYLf29U5sWdiBBkugPiuBZGb0mjC/Ljc++6CIYoxArEMpfriWCXQTTJS97Wg
BUwrFQ5GPxL2DDTzvjLiax9CIHjTWP3tXLQxLqnjpa6fQu5pSbSmZ7M+1LJDUWeM
gnqjcuQZx2/0EpiFeWU6zUl3BzPJ1/YCoNs42dGWiEXMqTyqScSqk2E+CfSk1yJ4
oUc8X+le5tub7ONpLDXuRn5qhlhvRZwXw0xjqU6xHCvQWbOzYQ2+P4SqDInFjAQu
JY6Yej1z6g/yhgS6dfyskUKGHC2rIAwhCSt8p2Xi517XBaxcybwphIkFjibIWc0I
hfuvHeggiQy5hA20CDHgK9ZGPtGoEvzpY54opQMpLO0ckIKw+f/aW1gwzNe40Cql
7JcwKYHPfOEZLeGapalQ5mfRKLy09VAtPumppa1kwX5+eE1qJl99eKF0joRLF9Ub
zXlUFp7IRahtpajN5GLzJDA5lBItLAs3Bnc7ZJGMA1c+nQOgsQ7Bj0NOXmShB49w
LNGme0eYczT7LzwG2DfsfTzAUeqbVJRXWEvC2Pl0wqzHD0XyTYFfUDb/3wwj9/30
o82KHXFC1QIYgpYCMRQylUfyKjJ1Gv3ML3trxZhTb4CSvL81zjlxeDsWBDe+SDLJ
tgoD1jbGEL9oe2Nr2S4fNh2jpVqyfblWY37nqHgJkShVNFJ1+hhjYP71aBhFH2Ik
pMDaiMtabRhAxfC3hs2WViO8wFBrFFNzRSaP8gKnxLZ7qtY5HaanehqoOyj4kkM7
OVbHh6rbkr8Xjlg1kAxM5eYXTTS4R/carJtmYhWs6wzXsscmcdcXoCerYFR+4VRJ
CsafJcoxG7RYecKrNzTlS3tlV2sBBDItp4OBey3e5KwHA7BNrsYbk5LvzYPj0FR6
e3kweMkpwD+HE6RE1asIaWPhsrVwEzKHVEXIpz8W9/+JL1OQwxZ7FND76rR37hSv
d5uCaZEKmwp47Sj+FIdGJhxZmKaPRdPXKgLArEFYoSu6lWWf8KpvKJJn08KE7owD
PRtkSa3GZqerpuKeO3yI7y6LoP3GDndrUcnSe74OZzN0iJ+6BZnxnVq2eW8CQUHt
mrrwB7GbGsrm/UDfx6XCoKwvRPIlTBShDZAhK8wZaR0VDlScfDtUoxIpVDZCz7fQ
LmRfZwO9Lkc7WuHayWIGZr7To6W6YJg3w8cuHJEhOJYLlHkWF0Qf0cSIXu+uoWI/
JsMPuocAskACBx64+gK/K/T5SR5Yk4H83EFtRv8TIRnAM8Q0PDUn/NG70LbVgzRB
tviVD1lTparprRimdAfFjl/YpUZ4ggJkZdy/238eGVUSZSlTBdZFoM3Q7M4zT2P0
XAk+/MpnT9Z/d4i1eHjQS4b8ZpHiOeon8SC3tLdTy8i6bd/cARRa1GCUWcQWt7SA
iI8S2su83emhzI5dEY0opUzzx0qHkID/bgh1NeHMvFZVXxmXtBnA6SxL+6htxL0v
YbNl91x/WVa2BJlbkSJFafL0ja3dYWNoyvYI7KNP04Vok60tRqgUok5J23UCXN4T
k7BbWPTAeDrkowsploIfitEPNLNPuIJdN9kWKvfGDPfhvUfyZg4RstinNo0vXhB1
r+lG90j2ZYHCEOJnaH//mGwCED9yzJGz4OAmqQ0wNykEvRnazZ/RW7q78TtVLmpC
y012p3IlgFIUxajGpoAlaf1izD9LcIQKr4XFD0/KkARPlr25vpmHf0U0y/blEwvL
aQ7zka5aVJU1g2Mk+6FTO7Acg1a1n5X0lg2Feue8Gl1rk+2KIa44O6eDfKkio2/x
39PZXx03oWIu7TEOJImhu8Vqrrq3TuPOz/Nis1rYvsRF5b3CzuFSQdubS6XxWcBX
xlsgiM6fkhbWwpikhHcFsj3+Tb3w+jWvUuLEkMnZfosajvPNjHTHE1IzFEYh67CC
TJsNKyFWVYyN731L0TPrvoiFzAr1takDsqwgSyOwPZjc1q7qovrNlERuPflLqznD
qg266DPV1xY4YuY+/3UTKsq4hf17J4xCOOWeqOIx71+E0ktyMwcDbgIaa5A03M5f
9CLCUv40vP1pNNbYoMij+DxFgoVT2L/rKw0tgOLYEvI9AsDAsRbCF/QSS87oVz4I
asxgJaNgFvyW2SDBeIsdTGu5k48VKK9/jPdt2BJS2qBOeLepSdGdM6vfuKgHMKsf
lW95AcdhcoaeLyz/sgtXx8ZtrIpviSGMrxk5JwO8mICl5dLhtk50EQVNkBaqiFPn
AbjmF2HW9MRB+fHloYDO8uJl2OslzTbzb8/f8Fkdv0GG7vUPQFoB6bkZspWnyv9T
Xjtw0w0TgH73l9W5BYil8P3wcRqe2XXozo5iPOFiDLL7YFtfak9a/DM2dgbqYJwD
mLke+AwX90yIten4GTdB7bYmjuCdF//Mrcw9YLUIX2JOlVKmFgc5JSNze2USdapp
jD1BAJA5+cQDgXJ3gW791+v9zHr1g6lHTXF79kICjKNsI6DCXcMKtRUOMuQxHd6W
nHpsHNplj14KiUxL+rhBMLukrGFlIESncMyR4GS2jF/Pe8Dobm1KjXAO8Zr4vTyz
XgYj8l1qJc9L9Ogmnc8HEtDnIIsBpHfuvL3mTLAX2ITmlzVSbxRq8vPf17cmCUYK
Coq1dW1DHxUj5jWQRr0fkvEeeRRUezUJaVAIK/5LTsEHg+8z75ZHa964RS0SYzvZ
QNfFxIGakr3jefMSB+KcOUL51zS8cHLOVoB6o8fShkHYjO8GQnCE2ShLv9/UrFo9
0gNDt/TBlmzDCq+IHFvqW3UIjS3C79DzcG75OEDy+LrmW5YGp48dNQB80wSJujFx
MYoec1sDR2AcDOnvabdzCHvEZTTEbDzjqwYMgAomoOLx5ghtzwVppzOCt4jq0UWX
ArNShlgc05VZTBjMKUWFmqzBdPkffhaU7i24MNE0IMW4w39y3xbuKcp5s3v5rw3p
522H9VAdkXBc5OOfTy95OgsmOgIvkQD1F+5OGHJjSz1mJFPNw2WIpEFAzJc9RvEh
RHYNJarTmjfgSWEImqSZfZKiSeA21N+P8k65YZbDy7eZ+DAcnhvB/vag/dZsaIvv
jyJuJKHJwuHDNv4+IJI+4MBqXrbKghZpLKj/Jht10qfRGJCm8VvLr7IQBdbB0lwd
eKAf9k99dGtwo+kVxpyYmTNzG++bxp5kPrAviSb+08VXq4YuO7aCSAHugt5ISXlU
cT2WxlWRL96ANEr2eTqUHX6VZNtxj+HI49nxo1iRniNz6g5WTiOZ5jz6RWpg+vJC
vpxCqIeq14eq/IFI5PsRV22oQ8fSBuw7BpDDjSW41+3FDtKhvtgeB12A9fnIgQ1+
l9iCYa24dolP2zDcw7Z7/EAVJlCLttPC0Nxmc37EAft9ZTBeIH27V1c+v+cI3vMZ
KL6bxeQjwgRZ2oyMSPLG1d49z905bUXjRm3NxHq4fUbt6cOkX9wZdC80JdfdhGaT
JdKbZr9PCaGCHVqSrzrBJkFBkOZ6eYLQKPCQL7MBQkB+PAOaygkpYTkdbbUV8Wf3
ZjTh+ke+IQKvpe1rrw7di0tUDN0uhuMtr0bItQBKUgzPs8mUAAxf+pDJ7Ircd3UW
YHHVUfzo/lgi4Spzl72t42PwfUMczqJctRUsLGsrMjQmtlBw7z9gc1KpFCKCAaso
rNHo6ngOsYCxUY7GZM49DFMNosOUw4nVI3W8bFB8gLSJ/6obwB7RJf6E83LH5IMB
GcQuwue3rPV78Govc8JwFe+eMl0h3y9kse5lgZ0gjbC2MwPu3FhrJg3gPOxAfb65
7IDAMmeddDZrSQ6ggsGLgpY8t7UXeaejyFz/IL4c5CBiD185CO8Y2C9b/Xu4imPG
EQrmCTWyuMEuJXZlK1u6nUg/++c+8fDsPDI3w7GtbLbfpgvZyDoEFSeLAiCe2kPA
SMeICFpSFTqvZI3PJyGOeZtbk0xAIUeBrrDo6jrldVYM3f2qv5JtD2Jk8hSuf5Zs
YCdBRT9LQ/t1dUlr2mhxbvSBV1CBDegOepVXbKmD8vog7yDG1vn9tevWX0UtC0KE
Gsd7Q3gndtHD6tipX0VsNUbM8v3nWu/XJuA4N7O05xKA0Ewi0Oyg/F179IKHx/SP
Ib5IN/UktnTwMm72vongt6ajbFv6EgNjLqFLaj0a9NU1mX+BwzCHQJddrXi+O8NV
wr6zv9u6SjAfAKuj8vX9Z3g/mCgiEns1hRfcFeuh5r8Qc4ScqjKK0111SQvnFBvR
xvnb9xJnu1F4/LCSMuOBFPwyhKHCoiioTM0Vz5peQ52BrlwcOvqr7xRjf7r86SVR
1l+y1TWdBAD4HTaohnF+2025i5hg/zFNhtfqA0CorIrCXCRi9XHUzQsSdtjg8jL4
I8BQzolehF9U6g94lJJAABQdaVU7aylwsvGH1L83vpWJuQ+IDArICWo6EZRvfqaT
4LhIPZ+jkqewBYywR5OJMoWl1ogTQgtqtlapcjNCMk7EHqIJwA+Q17LDdQl2NVjO
87p6wcIgrIgwKrIIGAGaOMN7En4fSAtFty0FiOBz8nZKYdm15fEZ4w+p7H0ccBZY
+cAnHmtDlmSvY9BdsyWolT64+r3KyFRulsHO4WEIq+g+I1ZVo/wMcBxoWpnrDW/6
+mGToXoczDOVYMXvg+rJ8QMNoW8ZhlpMPcn3Zifq/7Vg3bFCLHalW+AdJUMKzhI9
L8jJY4rG0N3nBrpLtqccfgtdzAaPAR66uKGCg4wIEVmhvJTpQrqElGqTJKvQEN2b
Xva6yJaWgiSqGVXkAoutpwivXK6nLvsprm/Of5NAbBXpe0GWRgmQjeRq6vhqWXP2
ThymFpPacq8C1hJmjTIF6Tu06GsJfHPozi0TYUHVhQ47CWJQCLIflZnZO+MfdmEy
TOwU6zW8zFjtefqbb4VPMt49u1sm9na7aU35PH4NipN0K+BZ/XzkLBU36ZZfStSW
ZL95DAjkZy2VDe3bZXYUrHtYdPIDwW5EDZcH8MtIAn9ZSd7HpRuW4lsl1eM+f07K
yQg3iZ24T88gYLXooQpelp7UFSda3dzNhrZimT2apC0q/U8BdaMAIoTWAEciwft3
zcV0KBcPx3J5kn6ayt/GNL7ySOH6poLCCVkaUW016va7Ul4m9DpNDiNQ1qO1SVhh
ehv9rPmH4o0NZBifM7h2H7Ku4JjEsIu4wWEEXmMo9pgWeFbbPod7Vai632Blbvj1
zgE9z9LVYNGpuuEf3g+eyUHzXPrzCoSJRCl5CcPuseB5xBdGdhMc8jMhR04exGC2
Jb6Jj6wK9k0sCgFr0U1Kbe2KHCW9ewG0Uoi+VKG/0voWPIB46fM/El2Ry0zU/gVR
5FUtvzFNaGm+DP4AxNsnSEagjKa3x9NaISMaguWyrvoHmKVU6UuoCkzlye+g/drW
5oRIZtpPApHTedpjSlp+NKV2j6w337c9acJ2h7SO4dr0uAqKdP9IyBqkpBAkXyVj
i5s34D9eVDnn0xjm4YCve8FjEkk4c80WrKbM2PPcX1dipFATF7KXXUwAdpUkVogC
OW8Uxe9c96pMuudHSXBVwAMeCFqljoHgq3ou3h77zAA3LGJdQYYOT3+nTgxK1pBG
+pqQRDWCKlakJRdt2CenKtEpRzUVgupijbdDhotLkWZ82aj+gEfawYBh7unS8Jko
FSih3Anf7AGbikKyGN60Ka/S3y8k8RUYmJESR1lEGIO3FNuLNBaTT78PNQeHoaSa
VAlljlVBHrOrSAfoRG+2pHMyNLdCUdKiMIL8Vcmd3oMaVg5wd8r6T7/si7XUmgQd
iqoAjmVKL9Pt532yg8TiISqXZEt+/OJ8NsMnOmztwdr3iDlS16dd5L3RFt7kzBXJ
JI49xfKOoTYwC5i+f8TFxzWacTTZ9NNwEAaxYd3QjqXyVWu3ogxkKK8nzU6YotdJ
aIh15fGmeaevgRQcBKGHHz6SeC5qsVzv4/8UnoHV+zh1s7xnJX+rW4y7KiZBlp8n
VmX418df/ALuh6iZsKF24oCr2FIwHoE2acRfqpIyu4SZBLeq+T1zsPSwGLaDsQ+Z
x3C3hnU0YstsBmITVyjNaDsICuQ6/6EHrDXuchUI0XTg7k7bXGzeCTK2XqUze44X
Dr/EHTwwtOqKQFOvmpu3JEP2LiX2mL0+TZTjhrTPeA5klW9LzORyZEEy6tG49SIv
sUwzIJljUwZ4GXVBKcnkVspLNu24V51Dpbw8kem847G7MvBJJvwa0dgpboRTVQA9
LES8NQO5ovirQAfwCHv9Vtf26Nc8WLNhpQXV8ICJI7bwzY2DzXFszSWU/dmNuH28
L3rI1OKjxM0gQ1QZWBEWgYqzsK28fnk25fjmCvT2NgwztxAsoqY/VQ3prEjuuQZ5
QvgDO8jVpRoiKCDHPnrjsRsK60t0qsOqPVvxQ0xxOayM3VjVE3ZJJl6BdPI8GGcv
OW3o4zXO4q5kt38dXiRjnyY9mA2Vs4iVPFj/i4ryWCyke1Pmw3QL10j9Sc4PqMgm
CefVNHhoRZXr27I/4S3N3LxWUB+EraINvuSBOF5gUUIkAndjdCHP2bLpmLqejct6
/19UWjyoX04P73C2HbZgwb6f2kf8U+h5AknquJR8ctufXyZmuvKQAUnmPGq2XkUq
RImGENe572ShqwlWiJiBQEFrUZVDvfs34P0nZJHyrbWBqEexkpTD0IziPtd0u7b/
UFX3g1ckTcT6lJiUsIR7SrafxX9LzMRvrQCVKLXbC2K2hA6LMXJtwpVa5S66geTu
0vO+fkDipMunEU77Wu8GpQKwi+chr89SQCZzLkICsE6zmVwOyVy/GC3XGzdJEXMq
WL7tUT1lUIRkekIvmEBRPFihQXb4h/fNvc/Pu2r2pt51hofVqmcyu0YKQ8yDzlZf
M+mbeLW2pXpyE9DVIvSj0oCKRK90RSJ+gK2Zc7GqIE53orFVXkW+D9qJ7Vv7Ymnd
h5SGxOxuqJ9mN9pBuv/Sd+TpIbLp7iYoGm+OR+rl9XaBChgutxtzJgCW1TRSPrOt
LX7UI75jiImdkRXE5jyMkj1QmfRBpTXhSpDwuUC1FmYnMO8BJwjgoBB9uDzxzQX7
LxMXw90l8A/8QloI5EncdhkyjdJdleaZcPEuqeVkkly5/9Uxc+sgDVOY81JEhDjP
5Ac0dDIjPMITk5CS+cIllxYiFVkHaov8g75mLndPis74NLva74s48luWg+WM54p9
jMTBK/SUa/fZAIeqnmuwv9JI4kldwEHou57g9NlYP2gtHMRUA7HOz0v5dzyvPQGT
2nifDWEIijfc/8HULpmw4W0nn46Ap0bfkQFGWQwNDOi1CLJZH0g9EZdiqiMsWmPP
1i2mk43MlJeumXAGuxmCF7bO3Jv89SQEZpeAamM13PufBC/qZDlVC7qYR+rVPosC
/FLBLE9Qwn3xA8JV7RKr4KmdEakJptiTch43Z/OxIalnNg+orrIgd2vzh6xOkqat
DjDzHgKMwgR9c9KEgrv2aLL+KEyokiOm0Plp5b3KaCRDJSVtZ5euRCpfCQdqwlhb
2pd93dK5J6ioMbR8ua5swizPRliDVaGX2pcZKUPYNmTYNoKmlxJBWs/ZNH7fPIY3
IG2Vn7vXM/EHiXGIwMpCFOYOx2cwmd75T5wN8nJapK0sH/+O2SgX5MNGydhNHmDq
tNbNUq6vJ2JAkkWGvTAppMtcS575YikjnlVe5lDsZgDUfVrH6x1g3uAzQTV84b3C
tGnrRwrlc9JKqHKlNr29ZP7AtnngzuwKr3RMbtsKHqfhpMT6ps/HFv7HQVtA1pOR
RD9aO0VW1ESSCUJ8NStKTbkQv4cL5ieIRBotQ9/vVBvol7X2Hhw/tdGkD3Icsydg
DjWPWqOJHp5edFSDXLSgJHLaScZL7YT03x7N7aC+W4qbuhi1t0/6BJUzHZ6Oym1P
JYKuFw/66RD2HKpUoudsGJRJP67DxJtjPjaLaJ79sDJ0pDgOG1E6AXI5l5i4iX3j
KltofQGeAsGe8+HY/ahYnM7nKePKB7azWyVF6b/UrxYjpI1XVJ9py9kv3+z0DAAw
2Dicpgrth/tJ5cHzP/wR8NHSDF0gv7wF/HtrTTIh7eYDAgvX6dZt3cqwkVTZcNy+
VdQtCa+fJYDFofC3oFsEkLDWTfga+6mZY4LPIq0r+HNm9g3tTfizJwp4zsEz8PHc
ZmPMJRI9NLrjZcceOKV9q9CS4/7RtZ1bWZvUyy1pOv3fSHA0xcxZVmVlrCqHAPrE
/jpHDQ/yD2nGw0xKq32BMfUOrcRVxjo91UVpcc9wiXN4GpzUc18Mdfaq8Riectwa
IHy+0snp8dMfweE50aI3nwuZ+QFQe7KX4wDJicEqrawaGGbWkzipZZuFp4FKv46v
7quAxfXGg4+hIlQtCszWqmEsRdQT0ISpa7/blKeJx0JJarcmsXhkZrI/p4b/hFu+
R8WbETETkbuWAo37FQLkzhvsDkiH8y54HqDvbEgoukn4mdRXY1BambkEl3vytb4n
Qzqv3e1xCNAkwmOwKAsDqvgSTZLWcRlgpjgDCNTfwoC8qyBSH47vdLdztfszpFAI
qQ5+eANJmyQguGYpKlwVPJYwNRB4qIkTACvg+h8gXRPzNLxJ9/GVoyLFz/gXRl+L
ces17vstDg4Nag8SnHjTXw3eHgT2GisIYf4m9iBp4piTfkxfGAp2JLZUzKPIoX1J
DtUErKRoI9ZbthmPqjUJrhdN/Kt33+pwWkqBbJKLi+qIvAty7NbX5YeJCWl8CkXW
57OM0pAyNUzk0AYQOb05m7AoyEC+0IP6WsaDM05mPuuOdlsp3vVGL59cBz+pbOi/
IFYZ4AleMe1SBkYQV7pmxq5gfa8re2fCbkg1I3lT5GtmZO7ij9xYx/BpduU+erJS
itAUI2/rUPeAqeaiRN+B9/QDJtPvcETExjGVDRIoHnv/SZ+dgamMlQb2Ddyf43sl
NVt2gurbljtYCx6VOmek9ZIdI17HXK+VBFiJEwxHp+GVXRYmDoRR3tkykUt4GrWn
XhC/y8vUcjP9N0GwmrWthbULbVKkx8kP4jbLx3xhOswiEPmNqWmjlPPd6SIK6oUB
ytKiq471pRn//6GiIorGW+h5iJsOeVe2zaxNgOQtvHx6JXcCfrYFbl2cht7suGzm
to66x8JIrhEN/tUCgFl97mwwjjF15xvza2BxpOvX+zONVL+DlPmdXXOKNcGZB0NV
OAyfSwZxjH3CJWqniCYUhyn7HyFBG5tLKtlMoNyUPKCc7KmlOWFVFEbl1C4t8eqx
w2veRXOGkGdYInEGjf9o3BCD3J7zDokhH7NjGRNqnF8v3SG5xb5ate7wwHizgy/q

//pragma protect end_data_block
//pragma protect digest_block
nfUxHSKzl2Nalc3q/bRg3NqXMls=
//pragma protect end_digest_block
//pragma protect end_protected
