//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TBMcKf1LyATFaPHsWNWPNQqa40yDdvGBVYAtZX4TXDovIecGZly/vzaIVeKWOhEA
5h93xr37/x+23MH374ys+5ik78lH4vEuK1Gl6kqAXUf4+auAfBPHtV3mGfpGOw+R
+R+7+sRs2YSIn3+mz+WQxjF9uWNarg03SAFxTtwKv84D8bNW/pblcA==
//pragma protect end_key_block
//pragma protect digest_block
PEW5ZPfoKTaTDtuAPtI712daIm8=
//pragma protect end_digest_block
//pragma protect data_block
aYPcOuz3nubPisamU5UQ6e3ktSDEFGAk0v3XN8n/djtZfmF8XVsxckEx1CG/2caz
sL4ePOz2AdZcis+Or84UaeSvjauXYytbhozqQkky0ij3nPty7Ed5wRmjVKsQwBRu
yL3XUxTjgD/rpVhBM/n1SbxQXjXLC+AgdeY41AfH+4xXPUDntbPliiGFIJIwQUd3
TGjwsQyFTUBN7Kfj+r/M9L7ZBE8VeBxgmykibYulX5xcbGuOkhzblxriX2FV0Che
lfhGEtfvAKfs01Fwe/W/T8p2gMrrYydf6y77OjbYj/sXyB4mdL5J3VBOhMqkNnrE
Kr7NSFRflwgysKLBEBElv4lDCPm0VI8kcb7oYqchTUv4ZNQLUEtDWLUEi1dQ57SA
B27gWNCHED9N5AjcZmPWDOkdmHN3j958qk6pxYzW9dguujKqB64JS90JkNuJLhin
Ofs15m/H83l39CQrQKqFyyGqdELJvlXgv+cotPWdwQF+xAP5VmnJOQ+XdATxTFEq
q7y1wNdXoOwlBEqjxEd3pNr47UFPibXnNzBpACigMVylk66Qh55tkYPfUsaSIllg
kY434WqK3+/AEaP7jxUj72LV3r9imCihfNYpmWxoU6uKia2vf4UNHz0QmbFA5dDS
PrV7EKV+/wbieWrHTcExHmfQs1HRszlbR3IJAb7pjOv1dl2V+bbY/kXZ8L06lshG
uTDiTKNlVdM7JNDzA9BvCTH2BFS7fa6sV0BHjPCwEdl2DBFoYgvv6kXhpYbKcp8H
DZp2OjvuCKgJAhOFI6idP1IWM6TBH8S9B5ZWwnaFErecS+6WIrvQ1gONkk0IfPqF
hKCbSXjioFShI0DCvQZfBAOBpbDVVfw9+qkKfnV1L04JcSwaWBGPSd4vk0E5me3i
e6aUmsY9ZW7bvQ13Y3qJnDo9SLjnyilRBIvH0AzeStlUpEDfgpd6Lze+OALvgHQ+
YUjFDnPXxpSgl/oUqCdE/S3nbwAQ45y29CYrPM7BAARhVl0QxT+u/xzXBZARc7GU
oaoB9z9F72pTWaeFoPPJp5PWkjup5vNHtiu4CcBKFQnvWst0ekkxk36qqrvoo0H5
fkrQmLrCfDdv1Ajj7RCrq+xi4A9hkZEvavKO/TuwWbv17Wiu9WT1d820X8vqqB4S
4o0ig7/HC3Sz75qv+EEBLomBm2T6ANWzWWO1/lZcqmUzP7/oQciltcUE9XMFywzw
jaLm5+FWLfRWbtabgprZvSWCth4tYTdSETyTwpTpoZvUUXkSllm60PcziiGSai/X
+tSRKwqrFO20QytG42pERJdflWtSlGX9dDbYxhR8yBUD4AsLjgVRbQw/us18ReCp
Lic/SwXEcr2EghROfWGnukzk4myTEe/Qh7T0bLI8CrcAdrm8/2hzibAnvVfl/QT4
YlXZWHWMXTcIKxqMsbvj4SeI4vL20Q7OlS8bxroVe4deVf6mjWyrHzHPAJpG3BgO
0clNJ/0AoTKbJy4d98QYX9PZRMSHSmkff9KyP8ZG71FxVkLNokY0QIa0N4s3vRkk
JRVYpdjcaz6R16IGzeSvUQKRf55TyU3pcFNSOx0c+1TAoRjIE0FCXCTCk17Bo0XO
HUsV9HQtPZq7JLyFvNV1JlHHKfAfXFKtsHGp275dsjKvHNhoe6t7ZVXpAwwZApBq
zR6Kgh9/rgm84bECsFFvtClgnVXoe5GAT3aVToU8aY8JAaeQl3bM/McsysU4rg4c
GQgE4EbSvmbEQwIpzoAqp0YM/dzH/2OJS8x0w132nTpujn4+S+TwvI/MMinMhs8b
KqnK2BV0Mx3E4o6/QHshb2F5lycpTHz4VMHWZLRiezlTyFI40MCKX5o3eZ8h8E/E
uAR/eWQnfDRHEehDiBoG9GDGDfTIX+GU00oGbz5yj2HzvY5boHcGC3jZ5MPmAazz
QNr2LRYH1vpW+iMrOA6f39lO+GwCti1bwNyi6NjxlbP11Tamy2FokHUeFJdIci24
KuiOswHB7bW8l5x9MdSuU6MOOmD/+jPgTS+CFJfOJiUQII0E1UOuZxiJM8vorik7
VcdeuA5OGMvDFCV9bu8LXE1wyUx/DYi14MvhNGvjIoxvew8D+8gIOSR5Dk6Z3v78
Bf9KXM9pxzY+FtV/Ai89bdq/QXUeLEeeZl6PdAgAbsYzf6RkzDsWFnlexP4j/5yj
L3KDB88txpUOERIDbaZk+KvXR2yr3CfYRO1UsMH8VufhUNxHXBLS2v1J/Q5IFmGi
ATTxoL1TJRH9iVuiUoEQy90ehY4DFcJ/O9IF2Zj6tElIAiwZzJsuTt13RaNUQrCC
N2rpl9dwCoRdduqO80M2u82r0jsR9mg2dHpA1v4H3gUNakmpixY87qdr/tRtoQmp
ME+pbqd1DgPxgzRDfjrxOQr3yZs7O12aw+51yJyP12k/prUonts76RpG2ITNe2FN
igYELb5FLsXgxAPx9aT8cXiS9DdgEWqAATGJBFJvBcQifQdoZdiLh68SpMIbOHk8
vXnyT/yP/PYBgkg8/8jg9nLuCbr1y7ag78suNrqAblZrVLuNOQBjuyX8fFTvJG0u
aTJUuZq7LoDavbBZMdC67v18q72DnHg4I03f14FaUURpJhNubMbcTCt03xHwQnxa
ltoW0/GBuBFEH3+KGUWBOtABp25H/0jtmlGEu7MAo1wNHu5C4yYjQEQir41QpHow
FFVv/wotWOyqSs8yxoa8m6nacm25ZEFeTVoARc7ggE9DbYMybngP3SzlTq+Q4pYv
tntVhXBzHYF98WihMGsSu2hqxoFwwon9RhR4ARMQyRwr1Xmuv4PZfKk3JbCUd1BZ
/oGzwNcXRQr31aznXOR+XnddngscpWACnSYhhULElqum86OD2bSSw+xRFAUj/H+b
nH3tT8v9dFa/tJsK+s9kSp+YcTfB2SVq9KsPiXix/1LAuqPybJl/jq8gdN/2mq9C
I3cfABQGD1e6SUYF7FbOgAJVD8grhFXoCxeU4Fzb/b5vC/DR5aRnK2IGHK6xx1o4
pnT5B1is1oMAXC6fKBY25mf32LfWUNi+M5UpeFEcXsgrd6yTc57XxkNKlhvaIrNK
aWn4nWpzJv0/YGIaRhHCrrKfrYI5NjwmCKz8QPomgNjLq2cabkMrzcoUv8T3YG7x
kYf3fLUpslrYV93RuQaLqLjg/QbkZpZNw0EAF1y1qo54a3TrMZ8vuhBAuZxdlVtB
w88FRO/RkJ3TaUXJaVvm7cpumRkuLyEWNoZ37xCJHnxvZalZPCFM8XXvF8eeRtqG
ZAoBzRy154nnLb05/KXPhEyvrgtaN3wBXkHeAdlDWgE+bnA21pHvKwfiyUnQEwoW
/ftllbWPohHfyGhLuidS3cBwEViAbUMCdSKJM3Ky6plEBSN6oQYpIl6NmpkuIA/S
2C9iKZmMfUPWSNFBYV7NE5Fh83373GNqwUwJQf0FZZ0tOV5ac+6EGnZ4JCIr6k8S
DwiKrRXol5Xy32sXMcATGzJ3aNPgeRv7gI9jdM0GyPLA4B/iBABnV1grZmH0033m
KOHPcixU+IENSRCKkbFuSf85b/xPq/QiTjwf/QSlrKmLY5XixPn8naK4Uitf4wt1
BkPrMLhn5I0bjW9Rh5hp3H6MGVDN/G6oqoaCj7upyc9K7FMlI+QITgDl+K9LcUXU
cmY1DaUosLynrYqnUVVYXHEEn1kkSXt7LI70hyQ8kXUm5s6pKVW0UhIwGeO3XGTs
zjmmHtzBbNvKurpE4acMMSV62e6wUy3FllnN/uBUOwchw18/gO6iIguLUUeh7KRl
wu3f3HfAEe7LXUJ4Stm4KrOIT6cv/0W0SQydNaQTIj6Av34iGo0sxs8mKrhTsxqO
UInIuPwm3eU/37WboQVnLEOlKkrZ1otSpnylaJFyaQ7+SLksvJv7x14q15DBQ/iy
pGd0ycJqyHxwtYabIjPQrmjZG8Gp3u1l3BLijh0WdXiwssVXkaiBv0hBb1Kpp2bO
FylHzskvLjQ8/sINj2XNWTfigeu3hM1wOiLOKbcRe1CwLGQyaLfVSpQGb5qkqTmF
jNuqvBoObFdeq/doQhTSI332RltDKJ2esZs7/F8BhZPzcNcpN1M/jeadu0UAdFPo
QT2XI6c001MoMN1v40zW/0Sxnlbo03+9WlymFawn8A3/fNQm9RBa62z/62IjGpJO
AOwXFGQ9JXPTxhc9/K3xSgdk/A+AIkdarfraHwHkWhlga4050pirojHnU1FWvOzU
e138NIusuRRIpLPrwvwn/5N2HYI3gJd/21xjHvV9lK0acH4IuClCZpnod6oqtLGh
zILeMFWD4/d0BB+XfV+VM1QkwydJDbhKihCPsmkf5kc1+RhrE5UriGxnSmVJV6FR
3ri33aRkIRZCysESwRqn7n8n44K6D1Lj7fzBuo62Iez29bI00DPFQJqkSSyretaD
/OxH6uYF+YWy+Pv22RfAgmNAGtXbO+jyY8CxskJ52oPUxov0e2/AQbsN/ZkRY+7i
3yN3u1oLMMzy5XNd5uBWsv5mp/ggSYQMkxpPBisHEeNVkuJkzUxpaxhFMNxgiAo4
52Uh8GsOw0RLON96H1dTHjhABnTYgq4kDbPMH65/8pCbKbcHdSXOHekJw4muwR8j
C5c49dSko4OLFt/nZExrZMbMAdzIHPdfP57j7d1ieydxmXgUG+I8j+RLV8JWRKnI
B8a+G8z6IWrlyuTwkUR2iRu4mqxsYmmdblXe5OTbzJOzOYGEnZeDdebXHclPN4MQ
89Brv2DG0EFdv37fQWgZwvmLWg8AQG4poq0noXkn3ZGVyMuqFT2WnRks3nM+2NgT
Zzb7a1M9F48MwAyhygbGQ7InD+jNCQaH16mJ5kBQPQRByNnw3GAXx5OAdQsYzmwv
UO78+Nuek815Jlu0+vn0IUuxgKPjtaJz+1vyOfOzD12mxp1i3PUl2iOSfpUdfysL
xeeoxcuOGU0yIJhqZSIQMkMHNukdBpfe+EEQgYuNepDDY+yNlJnm5+w7PL743niM
enLrZAOw61M/7PPrxRKMabXLcsNgY9esBt5ihO2OkDzj+nPg+C6EVqOAAJsPZ0XH
m1jNAL+rsBGy/yeIH8NyaQWgJAZWNipy5END664fRCl5JBQGW7IomZG3LGGSg5/b
2Xg0m5apaVCsZs8jvjdI3xvTG60g7ipZqO9Hr2qeeTCTdU3gosTSe8W80apoMOIZ
g1S8UB7um+hlTP8G0PP2FuD3s4JZnGHcEXstXpWejJ2LWeOqzq2D3IGhgxw8BUFO
qkVAQvgdjZNom8j4e1CLUdX7HYCkzx6Kr98A80P937VF15uP20QBboO6b6VvtRca
AZnRu97FLxYuJIzQG1vEV+ADTP04sMrVA15aszv4dfIDcnxlQ5VCtkwbbAU2l73b
N78gNHDsDWT6dag7nRhNqEXMk01IJkNejL+22jkPpiRGJWu+AkMDnPN7vhhronu5
tkuQxy6iDhIr8azoJ8S/w4coULnR/6UZbhMUQVob3nm5J+VxiDw8Zn5b2uI5MKm7
aHZBAVNucLct3GKRgk5Q8h17YPrElerrhX3lYcDGGHC8kFtTxfqiORg7blnSWRph
j0vCZCFqSTe+PV/c2WP5H2mtY07fgc72HpPEwvOJPPom/UhfIzIUa3UEijZsvte8
2T962hz+nVvo7bj2okSYPMUJy/Go10V3NbYop4rfq8IqB7sFnnGNuI6WiPr29bKX
By1xruZnMgBrgMP7iaL8hHPHUfhj8jqiXGADSVopg/lLGxIbuGefr77QFuM7ocXY
GJBd59TVM5N9b5R4JoHAZBKErTRqElz0nWYj8Yiah2L7C0RCsaV4YjQfVvrcOkKF
9P9lEc1Xpr/TMdN4R0wicb1FOT6fwGWoIZtIVM8fq8e+QJT/ByA9FQWcLUAK3Bfz
IdHd26FqQ3oEZ1KZP2eqOmzTaap69HyGKt5dgg/FplczgyoGKVxUx2qTDKGOpc9y
YoFVWE2w8RrOl+xkmWrhl67r4Hg3hBsly0x0n4vkeEJlboJ1tVvO20POoXf6bEhe
NEmikPD7JKahqVuA4MwP8jiSEPrho1CCOLJ9qWFRsz2r9j6zU4wfyVa/CFy1do/s
HXemVdtjemGLjKEC/7EiAYXTRVVQU0gcHuO8p4wJn+zncEHYU5SdNIp81/Ok8WxD
XF1JkphzzmpFePwRl+zdTPbhN3yI3lKNkIhtK1BwSF1hAI1nNHfYvBKsWwPCQsUS
ot3ZuSfVYOR7b/oSAcDsprYlws8kOHQGlU1s/R0XFRRKVViNtNd7tfbb9ccqsWr5
zgJKziuwpkQ40AhwAN60vbgwmNwteW1Xw1kWDZY61th+9MwoRMM8DcDX6Qy7S9ny
xag2cESuigP8/CZQVE1AAqf1zwknDcpvRHwJfPxSmnlxPtNcTAdDJTMvXGgz9olf
6abubkwRdZ9RUH2m1/xtbR5Sor6PNVTCC2m83ygq3WzJ90GCKCK3uqH802ZB0/dk
h8JTkrFALznLcZiB6y/PTTZ9mNario82YjGlbnW86NTrhwCB8KLpJa5oAIZQLpT5
TbZqgeYeHNbxG26ilaxA7Uf1dhnSnmWaqiRJxw7E36H6EMkwnGIo8Mf1jkTE5tQF
WkbUNHx3qetAi804MmRu+Ei5IWZR0sw17+fi1cNKbCfmGeMMnHgPx1LEnTI59L5s
Z1TEKTA/7bMSFgsCcglz7gtLBvwLgkBxDLrCMSftAPFC5qycjDyTmKHifIJaEPn7
eft4TVMUV8BDISQlSTOi/b9eNt9ET6KQjraD00qhIltzQ+5gzSfYQw4G1FKVHOzw
vZ19lTQlYqGbso9F75P9qCYqO4XfgObGyYTo4mj7rHvxH2ALJG2qi6drvAUdpDRE
bMXMlNDMHVh1DfSlWfCw4sTDuG/SE8HoUfG0WBlV83QKBiCzqZXCECdWPmBS8gx7
2ah/TFeSlAZ7sshZ31v0B47cK9m8uyQ53FEH8Ne+AEpPNwxlQW38SMh9NVdL2VF6
gyK8qIgw/khuDH7fo8JS2tH5q15cNqlEIQQjA74aIHFqbR1sFiv6Tb02tGcNAODu
rG7S1r2fDN9ARBYP3VbH4OZU9ip7YZxVIfVr57HaKOctiLRb9hZdmLHRwPdOdIp7
k5nTYk4mY/1nzIP+EOG+kHMEHI0BJc133xf6A2ZAgF/BJHSGxU6QC9phVwqZzV5r
rvbTCrEpCH206/BzaG7P34z8GOfwft+qBgIst2SCScrMrMlzyg7Wwb+iIYlfziuH
mRHHCZAsnIwrWw+KwLAe2m5oEf9lwGbAJwgqlzub8gy2+zihGWdL4oxj+nZAk1AU
U1nXBC4mTZNQb4tWtRjSSLfJayEN8AyUTQ7R78GHnabSKTWkOD5pTZQD6Tyz20cs
PBImxO4+Hh5+3pLNKh0EDMPqIavQYV7LPOAUp7QEjmdPfUeDTW2fAOIDhh8en0/M
FjzjR7GDnu3Ivi/vwAWYasGWgY1OTHT8CReiU4upOjBLef10ekkzbezVzT8ps1jc
NHhE+1kc9Y72g79SRLStTDFbmdeWSToqjG/xfIbwTmG9h3LScsEpdoyqNiSKVWY2
B/ueezJqQYm8j9tpLmaU88pLW6P+FQvWI1pClZrqWnQw0EZd9vfX0PT32zE+5q1M
o3ZCfdYxmJpWgcmaOUq3AgSjTuoa5crOiR4QGealn+dkZbkd2QcHJ+iv8RBVtwjY
RSVzWr2iZrxD7JuE+5nhmtSB/IpBye0D0anQpkv1U6WTrQsvzANhMji6AJHtXljI
7Br17qhX8N6ycAM1ClZSG1CtcGishuq0CJZw9dbkbIq15EZyHX4gHPp2QzxACVwj
mZuhlAEYwn2IceU+Ehzqcqv6t8eNjBGvTOv+CcLV5fccvtf1wHkOBNt+20PClLl6
xGYreW5QFiJfBkwliCZlcmNRTyo+OZjokRHIv5QcuxdYATF6HBoClmXgWIrFgPFs
TZrQauhuBohheKAhP99hGp8oVfMj/SEEsBvIFqzm5O0gYjRzn4uVfJgHn73DLtN+
VuTQOAsPj/AfZpmKZ5NBYovIUK2ePEN3m2ukNReZofoZghl3USKb+yIkGuEdQG/H
YeAnMpvUKx5FHg58zK6SbdHKAdG/94mHOWvpkh0y0/e8Ea5EVHAnDM11WbaqumBz
cosL//uHhQImJXPhTy+sVkvGutmMGZGM0dxedSi57BQA2UzQdM37DCDfK4OM3Q3x
2zKrpr51A3wDpNJnA6m7i/d0s7tfc91WoD0rtGqIPDcN3w/szVXT1yi9twssHGL8
n08xaU1ONxz4mrAETdcbBSyijS82jMOTS2zuZKmsaKAS/D64JH8qE0tB0rmlkSw0
stoBgqO4VOr7dws2lR/BUucAbw8yXGnlCd6iY7zIGhB4CkT1Z4syBfNZEguvGsiQ
Qu+15kc/YmLjXGY6uuCfqLfiTfrrytk8WgQQ97ypFoFk7kZO70MZ7fA6smidro3d
Izy84v4PGb2PidFWpBgctP/Uk34GFE/AyLwBp5Q9CzD26HdSa2sF08mSsnmy6+Oj
TfNABIoEp6mESs2hLY2tGOH/sWB9CqSZHAJ+BQ6CQ0d8+8bnYcqV5E9nZ/efmKET
xzf4RPh9+Bo0kSH6J527k6qrz3tjVVk8bA2s2HiY8fqjRjwIkAE+QnVlbyBRi1VK
vDy1fcbIpWgqPsBwqsPPXR0uEcg3mcxp4wAcn5LwlmyeMx4X96sZSlbG3CTp/lUA
Qq8/khrs5K6F1MG6ooCvQPpC0qaroSlVR43M3RlyHgWriYHx2Jq17tNoNYPzGfic
UVXSzMuvClz1EB0r4aNh7SDG0+55FaskolCxWxrgHgr+WK7OUDtUCnOrLts1Z6LR
/xujULteg6Z06pQ5kWuedzFHyzgH2TFK/Y4RVg82VhSNeZi3b1qqDK2D6FTdSTDn
Sx47tMQgmdjaNQ3dOZDXNzgKFlbI2F/O0pEBKAo7ItC7QMG6Mb3Qa9py6h/eVIED
/o1hCwut9ULiDA//ici9qAi+psAYtzsfwrNlkM51YoCfjbLBbbemJFfNtuFUS3Yn
QZxdwFLbV9brMJko9mzNmdmzJPLdbB6PQljaIAyF1+dik3wSZ8covh6z9k7+EK8D
Plu95ikydClJX88hbGP+aXxi6lTXB+3mEwMh/+Og3zrzf5eK/KVVRM3nEsQf4XuN
voPsAhRO7Uhkb7qQ3Z2G2rmebQBuJjiCoCCn7Oz8q8TKEun409rj7/BavdpVcFkr
eEQQwKn7X9p8XSQFudls1L+L7arH9sG9HecglmTk+ixDb/VKLQVdzbCgjqQCoSMM
DKFBhH/NZ9pVRvyL0tjfVbYw3xhnPN3zw+VHStx9YAHHfC2Sw39wsKtxluui+cAH
zZ1X5MX+PcEZKs/M0kinkEpJoYW5mPpV2cJyBbqbnFrMXPC/c0kxJ3BuetTDM1+Z
63a0kfpz9+k7KiAabO5YvnzpVMiP0aKju9K6ZV22xogZ5tQGjZGnQy8lftw1i56B
Y0pCYjl7FqUcRQw9YAQ/VR8xVae+hM19K/XXNYMbE49UPUId6M941iaYUu6tKft+
CPb4nkW1r/XaQZE1VcjBvB5jNlOVvBGmPlDgj/a2YQqeoX3t060uHfnNoJjL+fhg
ufaMDsauYwh1vYZg9sQggvnzJl7IGLmh9exV/f7QmuJ3sumrFc+X4CN419pUYIkr
u1b/nV+6HgvadJZXDsk/WDCL57D7//Bo5cmcA8LKB2kV4XZ/91f4KgxfX+U8kGd5
LFs7n09qCI/4cTIvuB1fyhjLceq2F1RlOsgGoQj7tByvDB2oosCyUKv2c/ZhQ2mf
GjQjG5ICeIyysI8+kJEkIjcfM+uStRxZ2cu6MyBCKXfaWnygnZFfrU97OuMhxmpG
XTUobt72CWDW90wEyOAQD87Y7GqtI4KW+qDodrxsH9hqRq60ib4WJRvuuDwq5Vjp
h7qv8NtfibML1qTMzvhqjQt3OUPdBU5bBmES9z3VGMkq59AGKOTNwlBPyh0UUxlt
AeQ6EAytZaAs2Ljmnp/DvaTWOsKO4sA0eJYh3Mpq28XOgZzatmgOmQ/WLdcafIYI
sJlaxZ8WVSGcQaoK19HZtT4dETqe1dcHqq7fdhsJ7fdspI1a1An1Kjy1Gol688Nw
QzBfVOBYfF3vTNVw5IQsRKm4aBLUnrXzdolCqCYmxrqc1L9sIe+s1P8Og22YtVga
7ZoYNeBskTWOObtPblUesLN4Rxj4ToBkhgC1TbJNR5mCFXlpnvIMSgV9/rDo2nuD
Q0Laa8jl1CJOPnyqXfIV0J/qFO5DkhtD8vrAlns5gWVHOKjjupi+4miL68DwTxEm
eTR9vxKpJo4wJWZTS7JpBollTyKtzyri2bb38wjfL8D6po4SaluhFfqojtApbPYe
pSzbKlDxOoOSrXJdpuQwr+AT44PrGHzsb81fkKjnWwyuLXAVToU4IeVMtyG5RE0+
uMeOIcxJ5jWZzrBPToFIqITcSDRwxil9W6KRLKLnYnlWoY+yFR+me5opP+CRIyVS
mgyys7h+R2WmFanD4/zziglY+6/OAFg7y4/uTxs5OjSnMfGVDWGgEd6PBOSaADOw
p/eAS12dDg5Z/iSmCa8y4PGooF3XDgjdLMPLioofPuCtK5G9USALydKmE2wO6SkW
T6WB8yyGAmKbwUX/e87kQEveK2pWKAn4PKhtcwDR0dUal9ck6tCQ65MdxwvQwH+a
3SRlBdl6ZzwDMvKbIfd7Cw5+9ayCteF/Sqxc9/hFakgDnz5rm60QchmnBKgZYC3X
m4AxYCZSIO4u5n3qgkIfBYWg1DMFKH4CpSSLXqukC+dxS59QiLolwlK+o35c6mqk
Er7dkPHlT1vzJwRbadZ8uKnIx5Pf+LyHadP5iJwmtEWXV2hOV/IXj9JAzzoO2RGQ
QhSXuGDl21LGPyEqluFlhnlWL6FL2CYq/LA13TrzeME0Pl7uvixq8seB/IPKlxxT
rJPtKyh38KBkjs6eZuZmsQn1MVCjrykRQb31n++/F1etLGn6obHQtPmN0p7WQO/V
ZbuqlfLO2xxzy5a2ffd3S8YDAz2oR9bPCQ2Ys5j0aLbBVvwS85wk3gXVG4Tqfhp1
RdvnbAakyZOC7LM/5rQw3Fj0SeheIhSCv+9vVvszI48xNJNS9nd2Kcj0sX8u/p/v
4sKtWaXVR+jRLHpFpUb/n0LU3cSTzWa9cD+mzLRIw5jcEpjrOitEmrWhKJQfAo+O
O40xrRK4A9sjCk+RaWgQZte/u2s/fV+aJkCEnAnhmkamZls9lAOVmeySCmY5Jyy3
KKRTsicTf7P1ADAtMNA4gk7oXSLuwaRSicS5Jz3H7ip9ydop0BKG1magoZh/32ch
s57shddgD8KFun3uYCc7eOffz6d/2kJXodBpnpjUQeC8BNvihY5qK4PwTc0E7R8F
NlFje5t4coqJzWIMPBplT7WJVFiBVCct1GiToETGdEHc4KI2D81LZv5P2FfnIxBy
C2IL3CFyrQi8FdE/IPTS+lewV0uOPVU+oHyJmgOZ4tHPLramb1p0dkUe9xYMHKwC
i+ROr0++tya6c0zP6Vp5T38u4w2cEzJ38Z8YAfYfmuaiMTFv/dvEjF0i5jbb28OO
31yY41/IGbDOT/Agv1R+F7s+PsHhbrD+RmcTbz2E+1Fn0GvwRyuR8BmrNW5xrePX
7wh7HEu6NRbkBG+SU23OrV8OMXPOAtSIbUK3vGOHco7s46fE87OcKeYNIVGi89+c
wkeC3Rvmao1YPh+S1BkJXtgObAl4mUMkjb2Qd1dZkrLHUUccfKbiybCpMsQ5O+2i
6QwNvqkMw768YlC++g3VbIYQR7+io3+O1xUYCFasVAWkHaeHqLQ4Eu9xzeOCoVhD
pFv/T3TOVrd4BLg/bndoozMCzo1noBDW/y9aRehfT4vaeZVvDeOFACmp7Olhp+gS
5y7yChg9rgwqD0e3MtXs9+9nT0VMhT7jHAxF3KhCTCOmla/h4Vx95sy4SDLYrKRk
vTbdyKoVgUZZrRNQN7ppVUy5I812IF6Gc/2c0bToN6F1ZjXEYWhqb8KwcBtOoRMq
TeVKDWttwxoQfovKVWl+OtixtN+SjoGgGJVVBgAywM8gKUI1xe4gORd6psxJm2AR
H3lcC/My4gNZxdYn5y/fgG4agTfgd8Ws5iakVdkGJ0pHLVmjElbPChh9EYdQw0k1
Jwn8zU27C/GbeGtjHE+dtCUHqRH0ciKBIqUcS1XntOxtENQMz863Swdi94RwXVSD
6IIam+8NSgHTHmqibSKHqhSKhO9yWUPrzdkZfY4iSwSln2fHa01jydMqEC1FZStM
OsasHNZWBAR1HWTUQoyOTpndorEOeYqcPeGhQt9FMWRA3U4xO/6Ft0MwCVySonZ7
dOtwAwcHTq7x9GZJdWXlbVcf/VLv4p4RZUwnpjFvj4SG0cKH2dSxp4psLYry2fw/
LPyXQd3FhCZzL9A4UNdkjYMD0PQJsNGkMzJk1ofWIIQweVtMiEv4X7HDYOR37qLM
I3lXxTwHLDThH/+e8uDiQAvk9tUJPDUgDyV+qDtHytdmLksYoYYBEkDeZFWgV9Sq
CW7FWkJ5BqOCZz+N6cK2KGuc2m2mVc3XJd0FFx+XINxiRxKzkFt5m1LwKW/XG4Wg
1Uo0CEUoX3VizbXG7KffabD1cb9GGkajwFPbNEvqLSE5EI+ZOyXJoSsNDqyKJaoI
lS97NjA8SL/CkKsZCNX8ZlmJcNbxlp+OCduQXuneK1815OgzOjvw+VQRLI6FvGBW
cQzzPVoBNNk7Ah3HxntkXr6iqiQ4S8tt8KNrhnTqQJmVS1NsKtDvR1qv7bQX8rJ2
sbKf707YC7tLLhkC1WKIw1dz+u7vRN/L/BkRB6Apf/IhLolrUCKqWrEM5Yd8zlrV
BKk5yITOq3RhyjrUJIJkXbf6UUYegdJgtu6z0ZnMQrpXaD+lPXMYHDKFNhPqH7vC
rNNGP9SpqV5gcNekFVoycHqKWpOne2s+vCi/EvoGPez+K0eD1t9bwmf6jo96wwhg
cPgIvQ+gJmQkG7r0TO2n0svJeS7Fn8Su6KHfdKNYi+rQTAWxL1HYThTiNAWETYFa
nWS2+ipBacsSyBHA9l/oVu/ryQ0X0O3fIvjZgAx3U6aC6J1DR+1OwesT76Ky4lbF
nyY2pgvYRoflzU2GbGfKCJjimgItGXB0sxe1RjyLjg1XKYRnkh4+4EPKP3c61y8I
5fQ06xwDVAOAzTRTTPuaIAc8t8QEv6op1/iqAJGq3scPJZomtpE1Ulx15w6X+22U
oP0aiaNq7gfv/anfER7FJPJDpbw9ULYLNRQsO4yMF0Qmapc7qN+/Gfgwuwi8DLQT
vvUhdFW6oTzkJPrLrULSoZ2fc/n3iAqMOzLUDyIkYyxjJcHFQEf4gUTYleihCy0s
pP8OtMK9eDp7GU9duWT8ulDCAnEW1F+p3tW+BIqGjsEIeMaVq03KIcjz1mQnFaCt
kBTGtN4lgUoIT6i5h1SD8RMU33GKR4rJqcJ1t2tCtx7yxTiJmOCEOWBC+tBi3Ine
oCeD3K9Ok4/KThPEkJk9Xd+PpTDV1QpAeriN65OJn2DKp3iNvxLDjhA3CLfCycnt
fdQpILGhJOUQtqy2V9tMF3Dk4kgkz1ahstonq+GWGPEoQA26hdgDUXvAuCrcaSpa
Ca1fmM2ZIZQccImZHV4ZqnWv+OJFT/gY5gGDwfvpWeiiCuUfAULxQMlCrs2Hau5L
nLTeE/tZ7O5apgwzDwOZ6vTtKQpHMiCFuLa61xpKceETUzo6z9UHKGpxBtmqv7Eu
Hb0zO3JSJ3gJY+AnC93JHblWyA/hBs6Nn1KYSUZcVz94dteXt2a7A1w8TGIIW5Er
S1aTvhHNzs7wERs2sL7YovciUL0DQF76TlvU5GNckm1O4U4mzPoUBSUD9cu+GMWg
GKjX9FvApfTzoaAbnGU8HlQZ0VevRntkx75MnXVMi4LnRNGyxIOGehu1WEhpNtUK
Hl79JiVPNn2F4RwOQom9xVF97KXAIrDe7Ikd3VYxyBdQV4PRDuad7PVAJTGbYw8I
kS2ZxF+GW1scHpS6p15B4+yvTxxEE+FMOfwa49gc/It9XFnmlhZ2j1BWtqZY+HQl
R01uZgc++g8znERU2+ueBQjsmlfIm8NQycb6dTsvf6q28JphDQFaTFtqM47O7i2u
FIMbHvD5ZVpyN394mHo1i48BwoM3drXBpkY0VyenUXFxPUrt9PNFFWKlonh84+5+
H84jDPj0t7X6bgNvwF91Gr9Lu5OBROkEThxfUgb1zOHduNV64w3z4epgAQe5Vx/m
sP3K3Cidr8yXm0YwhvyDuH4x55DE4vy5pdF2b7ZR2pDMCDUVfD4JkQMNqN63Cfw4
0UafB5KYtutcLZl+L3TzfkRXvDciWEt37ekDUlCgpJXIqVPNGHm4pX+HCURR9LGm
yjRqnScQbNpxTCnb+tgNDRrcAqTP8A82oSsoBhEx/SpbmZ16kOF19G6wIK8grOGo
9MrKUIJzpoNRnYuaqtj0ZJFk980jhKOiyOEjY3K9oKafAoNVM1yTx3qOGt+zua1U
R4VxcjpPiDItMrg66MjX5dj1JPF4ONq7wTI2yBmvAN5RPTPCJtcnvU7wP+o6Icdq
a9f1daVEzmZ5r0BRBHLfcfuNRcRbY8qKPewY/JWJsq1vZawbK44yq07wVKwu9RI8
qykSjg2FKl9cmqb83BV2iF+daLNh4Bvq3fp2wnlO/j8gTpWs0Z4qm6pB4Tc7ZUgg
oyoTJbcKhxT+HpXB0uCdPR39W1z5PcRs7x47mB+Ne+poXrXd8ZzhRL5vN5DU35Mz
h5KuigDjAW8kMlWIqzV4MCMn2oagDABU5A9vkWlEpvWoY0qoNzlv1IhMvjvJgJYY
f81FFT5NKI3F+jp6EbvtzOjRdujoxYLnnb7gDrB+zNVy3DSAKF9jKHUXQdefXpt0
dzsVN0Y2KteLwKj4EG3X2FTAZefBjegSBoz7b22zLS5jGS8FJV4LTA6UHxgDi/Un
4CNQ5LfMpjfvD9md3PyD1tkg1Q7bEsuramx6RpVxsRBqiDqFq4wP5whKVa3/n3Tm
BYwuaIqJ6XYH8pqJeT1vR8OiNRVfYWzoEJtMPqXZ5Y+12wqQl8i6Wdpbv/1/gpji
lfL0a7qV6g9D/HTLF6bin0+jFYCZXxR44Fe6qcRES62+RIDPE6PSLC1PWIiSJ7WQ
AdD4JVikmFPUYZ23HKKbyfmvqtwhOCChzuxQ7H3vRSDoK5XnvilTylvnco9c1uUy
80CTJQqbgF5Q9qkBXp0OOOwmzPVw1/RcAq3ETxX7a2zWifs/Z5Clk4gSlIMEQIZs
Tkl0q8l8dNMMsklrBxu6US7tDtuogBNl8g9Wxs/zgZDgAIXTQtQlfhwrubRvsI9Y
Oqli5LIbSwtHXpYtP+ssvbzP3ZNGmCLI5ArD1Xbqumd7ppT6VG4Q1wRn29jeAdJo
WNRaH5ma5mGPJUHCYsPK4f9OlwLdF8gnQM+LlegYwhD65nGbop68iVcpkNQAzdW3
5Id1o6xaLEuLpu2J0pUIgFt7mB9VmFVUTwZAWY4C6BRQafZcO8j3qWmlGcFcufNy
JPl0HkbfbFIWV+fGvro3j/Lkfht1LHp0TQo9ae4F5U5mILrQy6JKf29Z/Dsh7BGe
DUyznCH85mYZRqmRF89Pq9rEeg6kUuQVeDIDTvzF2QVVernivz4OdF8SDRgJhRb1
jUjas2WfXzMkJwAHeZb/9JusOjExaDhIKCdWNLEFfbwD4oH/uzXy1l3xaf27zFkt
qz1ya4VrptYSmVayJWRHUm4gywS5blnXWfX/ddRPO9tSjTWBWNuJ2kAG0rdPP7RX
0RX7z+BIaUx88Hk44CJg6MftpU/F/shGByIelMM6WsIpiPPcl4W7qf43lh8hYWWa
xAo82lwCwE3cFBXTigPZ1+D57KlxNibOuFH8j6IlAvWeOPuFc86bgqQXpfpPmpNF
mizlamQpzYlpkQjrO+pyMsRvTxndafR50obPDFdMpsqn4pquACv8Yi5aXfkBItcH
MoUG6Bm12AzI4hcIgjbThRLTn8KluQ/m4PtSCvPWFKD65HPIkFpeTV2jG2c6OuDf
Kck3C5BE1qRrv3SPeIl7qbYNafWq1+lgGRswp9zyihNAXi0TdLQuCfvHeMjN6KHx
eggamwFBP6Ormhj7gp5jXXHK12LNgflycp1zKF8SC4fMRUJvzNaAPLYposgCplAe
OzrrWl4SztNxhg4rNJvOqKgZWJw7YTs6ofQ3DVgOrsPQbbiN8RsKe7zk4cO12VpT
u9TDHTFt/6iaH9K0l5pteZuwV0phK/drTyLJVMbBlQoS1bf+pfv5jxjK1Qdvz18D
Lq44EU5lWP9j6b9SxIY1UpgYFvHd8PW+SSTIqvASbnuGwGEJEvbcK7Oa9uqq/btf
IDWKTaie7QNZ2rWUIos01WFeNyp8HcegYZjvFcQHLiodzJQrlwu9DLWw+KRsoY57
yeQFNhpOl/lSwXhLrzr/q4FTLDdhyx1KlBCLPfB2W/wCOelI82cLcJP1kgDFoRdr
RCScISuPSdX3WTJNcSRk20IKO8nyj0z8+qUwJsxtzhE6HTBzM740wyRoSuZbkhYK
2Kxg5acOYKarmj6/IVIYkRL3xha4QXorR/XvvMqheSl78RQydo8zJIRiNXdq71Ec
e/5n5Lrfa9fJyLZtKygf6XuS0GsMfqTCtLCTtNfNSajDycEfNLg+tsWkkbDA03h+
b1vmqt45+yC0Gan+uD8SF8vL5FBlI8QNjjZ0bCa/3KCaeHHVV+nsPOBcuEz235+J
evVl+MUxAlqbbrHwhGC6Q4znB0sJGTwacVfvM8cdatDN4Wmf0z2bwZJXTX0kut4u
x4PruARmZ5VJ9PGOrnnhQiOKhZMXSS6/MP6thIuqWwNYnRsiVqjb1PqRMj30zSef
wPTB2qwCfFAnZn9BekjyAmf5qi/Ikzti5iDctk3puOBcdDYWApJ5AIjOd0XNtSYA
S5E/jVVt/E8yMCK0H9h3GgGuxUtWRjoS6nEXojFPVZF+OvryMTofs2ppZLCQjPtn
JJ5yVDz1Zqpx3eNLVEQXpk1kiSoX7qw0AxbzqdjyDYYiZ7Vl5yve5oJ1UY5M/epS
vVqumZ1DYVYVqM3loUD199URWA7j4eeFSQpm/1BA9VOSRze5++sneCEY44+oPr2R
ZzpGuawph2fguNNSuL0vZ2rNx4Q5gvwSR8l4qMO3qsPbpr/gQYe0sX5Fhi/aIjVQ
80pTsEkjQDqJpY3YNBpcz1ZW1JxGyRSFWcr1Y3AVKDXYpmgs7yOeremmZjnUCW0o
Z00HSkT/d/tAfVKETH6+o+rXSNlXJNdvdUCSWVQqeOxsxIfQMc918NRsJWw7rioX
jgr8qEpW+WoXXiy3F3wTzQVd8ZJUvlwpzPzLyb0uy0OK2eK28KIBovj4Z+XhWkrV
xlPLJtBzvENk0W7eTqcFiaE9Evtv6Gx8CB/1FXW7R5X9NaDFrYtZRIYu58cBKh95
1ymcF57LiP+XyCfWXC/1dAopeSoA21hx6d8P5525n6QGDdAEU5iEbbY/qlzZAPpa
GFUOGmPk3uRc5hN88INfqTiE1M4/P6vara2gFaImekJ0TYDZwcQNEWQguOriPw47
yFMLSGpgEtXFzcjjyShf8vOm3E38KuFSIC38I7unp/T60U80ZFu6l5KEedVG7L+G
6dGNEe99yF1f9/LLECVwJLHvkxyca3SRZFlw6diYd3rLneiGOKrOd5tDBoN5XLaS
OyGHAWnJskExeMv3w5iB1z7CAHrSUYM7tAR25xv4mmW2w6zD+e7oFsd7kNvE1SDa
uaR+pKFIavnyQCOMF73jovRKO0HJx9PoJP3nIkIbWpZAmXEJgwtkTQ7R50nDaC2y
qG9bdddZ2F8+e/vZX+w/mWRNU9rzRftaKdnTojs02BkqYYivkVmXmt7EIAXNr8bX
zFmNzkgYyqQdTx1RqvTAHUheTrizFJsvWqG9gO19D1jXC65+5mT9+e48lqpCrole
w9uoXS99WtBGNOheZA3eEcAjUsfpfTiM02boXKrQ3LoDsAOlMn9osJV4EFdf0RfD
joVI0fQzFM8Y1Ual4eUX2T2UZcfkbfnsE/XGFxiUYrHrol26nDjNXEdyuUmvQLIe
wfoBHxVwC9KeAfR5GLwQRV4NPqanUlfpHX0PX7+DllK7xVrAG8U2uo8kv6i+Bn3X
P7F7wMSI0q3exJZfK94yTTTeAEM0v4QXQJT0ydAfC4uKeTkanAt6+WbIkw2TjDTz
KpV54M+BohhFMzEkwXm8queSXXea+Nl2MJhiDatmV7iCi2Z+oGBWRNkbeo/E0sez
9BlzXl7WUqwXK9xi0Pv49cYD3M5NpEGbT6m3uF50f8r0/na/mnkbh07BVyXUAvV0
2HOeoSKlteYLB0ZeRr1ZEUT3BeQUA7QPSA6vj9Vf9BP+mrXPqBhIFKGZu6B4s7r+
q/zlnIgqD6sQfG6Mc5zRDswzw4eQow8mJRhIiPUneXEhCH5U637uM5Rk1o8qpJ7J
2aSinf8wI+v7gmN1fzziatFLLN94zbA6j/aBVtk+fCfz4mtmrN33lVXHMvz3qUhq
I84J9M5czVX6FS4IlRkO1eZwS5g4jW/+v6Sdxkv/SKqCM0cuLpAWwhim1IJwBmKo
xadimqsd9C44fTnD4ZjSAuqLrZpK7hdczDttd+Z+PPRuzlTWo3/B75XCSXFsmGSU
ZFICa2zjp9bR3sFnP+BwEN6+iEIQd3+M5yKisMYMkRlhe3B8MCR7PKWAuXB/TS9X
dZVtPlfsFF5CX6k/Qc+VV1trEiGMF3JlalVEH3A9RZi4mO90691g3SZDINcGWQy5
vPHPUumpA0AlkZJM74fpNSlDTaoCnyWPLDL+uFgNWwtIpbyIGcJhtQS+JAEwpzfT
VYkf5D2iNH9O/349UU/Y5qQUoVTSYQWSmSD6RgWqu0iLj1ieeFQxD3JE7XBv4cui
dJ3cDZamtJVCreu0n7IILy8dfWFg5tMiGJCanPi+TwqNDE+X3msrkf405FX1baR1
5F+Cluo8fVFCRGrhtaI81j3qld6IJQlGyszHbJvcPQ0Z6bx29YOi+xRPw4CpLUZJ
ssKkwuF7J7J8hObdPPXGn5qlJQp9ytE1sjIzRwpZyy/Mw/mgZH2sjnW50xm2bM/Z
1w8+LCBDyUwPKEQPdeJLd32rkLij2/DvffbjNie0cTxQJ38Fgt4Wex1kuSxUj38M
TYW56GZ3hXbS+wjoN0LRwBgm1zv7gObbmyLr2jaWz+vyqCG+DTV8Ob+JdaUXlNzK
sTep9C+N5wTkilOC09c4SjqkqR63S4bPNt8aaJLE42oz0e1QsSv+cU7h439KCrjU
D36OYhT/RaIxAm3+axparbmZrAgeF19+MCO6TXuihN3LkDmGa7Gt6mC3wGmMvgu3
seKT1icuM06GBGNGgcQisZlSjD8PJQFopPMoDD+R2J+iFdRApf2m+3qoYWzZ3Sjw
bnJSuBfcGnIJi4EfossN03IDhK2R7yqaLM/mXhIEmYpjaf0NDiM+UBMP54t4C4yS
pZB86pc1utigM2kh3oRlT+DwSem5IGCpTmKRP2TCwK6rQ63LSSx4YRDyezc97bti
r6W/ajdL5JNYSboSKgAlo+Gli9/wiQCDITeHcwrkgXkz16i0lPaL0VHPuTKqFJ32
FfIg1OTJSqqpVl7LbMLFGO8s6nX/JjRTgGDbMT9AML2DBiLW/wYy7XUq+Xw7VTco
IpJesBFwAxjhqJyAGFq1OsDzzS6p9yeahlxJN7aBsGQQKR6D7oiguaAH8c6Xdisv
cYVJ4DWw8AoYdlSbZUS0mrSErV4J9W4phJASSYn5gTxMvzbfAGDGMyQIkW4X0gPO
il88+Wx/tbVh2tqn6n6Y8vjsnzc9h96XdBMgHwn01O/oCEKSA1rxicIHpDPMMnsM
gk/oyhWsV5BjNtBkQniaLMqAgI4dfcRqRzvri6tGlJPraGhoPRjHWLNow/UcFihA
s078JpqLzUf8JiPTYE6WPxQQaNJ2LBfMwBQ8sEXJN1tN/W9y21yY0pejaXMY+fXy
9rh3jr8AkgWr+LBiATuXeXMYZrNSkLWCtJQL0ifWa3FM+HJmYOGsgKWDlpq6NKUh
xMn9SMmHqrtPbqpTBGVchJsALpclk8wSDhuuGnC0HmDXCZPhc1Pn6x7jm/IuVfXH
TTcRvIOwMZvBqg5cE+pBN7WdQnxfQoxY7BKP0vMe7kHG1F70bkyOqALyDcIEfyf/
S25cpltTJ6W1N9qgHnsg+cBFVCy20w7jK9NpBJmzBn29EiF+4EGrNAnI+NYlsR9H
n7cD8C7QrMjZvoRyt7WH01KDK9lmKYb6Q0JWycODcF0SbRe7YK0pmF9OsdEl7Dr2
LKiN7aDpfLGIaOt0mCPfQ47f9t1GGc7/GpQG4xf62Wg3frAOflF2L7/V8vEjHkGs
YCM8bDKjSQ/3jyqJEmdyiTtxn0Hn5fy0Cwq7bCjh31lQx2x2PSBaXyjgJtmmmfUO
UVX00rumopp1bS5M5hbCftvoeVSXlBWExpuzf2/9jLr6U+xfR+N2IFP7NbNsYFe3
bt79uD7r3jqkjACXHkmDuDPs1Bf6CB/UD1aABD4TrXzVlYFNq0G99XTqb5Om92ys
nPmvhV8hTEBtLa+2e+LjdPFyZzDl5pT4y6K1CHw1ZqI8TpwL2zvGYZVTeD4e7ah3
tWZD32T8y2suBQzbuibxoj8BA4MoNEwcNAojq1mu8Li0iYkN7HwvhVwvm1Yg9S7m
IC1QK+PQ97v57BOw4BTKBGcmTrxdMC7zyTC9IwLgTX3G1gNSgQQi/4HVaEhFohAH
7tYUjMVhkNrQOGdZAnXw1h3gAEN6mVhdfVXpNtG3i3Mel2pyv+VI8WfrKW58LUcb
jnPa8CAcEnQz2//qxTsFiIKKchX5hEuSbUpwwxxDAiUAD52txxASxGhD/VAR3CFZ
/9nDoftHcLlHjlRA8VRdYUgUzaDHZy8OuvyaCcDlezBq/gTEbsngZOJYl0IZqCE+
15r1LlNMiXcKsqYxtTIMCvF/49lJsOxhGgwuYKusZ4g7U2bA9HirRHeWqaPoppwG
Xts7Y3kdBdn/J0lPIulpYXF85sW9IN/kBRdT1N3iea4TgdnXFxSucvzs7HtbYc/K
zIEouQE+N/CsgGEemPDOxWXTvZqksUYDHD31WdgSNAlLQewwIv/dwvrGf+/44FXC
3jnxPDcIi0CZpOfAUXgwVNGbcKWvFYPJx9cA4mHakGSqC7kdprMv1rURFR4njpRe
kQcoRGeJwV/HrMPZ1XVK0N1mxaUpgJcwQYmbDNID8d4/z4QszoPJcuYZmkIPvE7b
jb8nazh1iO9l3m/42l4TODmVyXj3uPMkRXeLih/DiBWnYAEG2sWWD6ZRZ8w2qYAg
BhV0XCSE53CTrXDI/eaQRDcScVnlEiD951w7jnvsEFD/WZ1ufR8wgFPiRMqBlz3S
z3Hrf7ZNdHdOIel59NjOJUajI0iQlj/kBBKnxCOswbMlYEz3pDkl/NfhHZUSdpW3
2BYCFRlU4EFpSW9iFW9VMc3XmscvOdAL1OToqaP/L6mlcT8u5c/r2mojkIEtIQDt
wltnhCSpnQis78+iLOYE1tOX0CJ0pMfM1wWsz/eXSeEq7EfD79PLIQQ3ONuoh7tR
0LESg5Pq2vJGVztpVLJBdPXXXbiMqUDqclS1RmCq3xztbSha/elRQpcXLwYNpA2N
zsq/35uPjGVChJd2HvLM58MBVk2TEBWNiUVBfWIKo6iO8ktL4qWItMYXnSmnIR+3
qdGiK+R0IWTie6/AdGeXQMs30e/cUq739Uhx1pEf6Q/V2dVGgBiiqZChzcSOg4+7
/Xm6xgA+QoiAwP0YZVAMhR5Ph+tbL/gCvPezj6AYJD61nzF6Cfgl9m+Qi22WVxcy
bLEOFVY0NKuQsmt4FCmBVwRXIFDsurgknLbvJBpUobN2ZNGDk7aUBoPPbsSMZvxp
tgeqUL5Bet2hcpLwjIsHgek6E7q42vDdNxBtsFWHaFE/+pWCnsXIFy34b+6TWVBK
Z3U1Vz3vI5AeKIr3xL0S54yxV8ztEY4fJoA4RyCflH8TKhHQzw/s9FQHhDgCJuMk
m9bN4jk2fcoXXLgN476nBsqjIHxzKp6lmhcHsVMB8hXOBBy4zwvaKQSObZqWB1Z2
+HGg/xSaPY+kBxiUakmNhegSoutSZeuEKLX9zsj1U3X7v0MXqS2X5QjH0Bka94m9
cXQgEBFv6jNbWPt30ozm5jf6HY7CgpKiR+AhvLhzW24o570pxVXTae7ycn3LFjO7
PgMV2kmMPpFjmmhOg/hizXihnED5Ddcg6CDDzqeSQFTe+gc8ErtOFzvU8H4W0wZb
7npRemCTBCcClZHiBiHUVaTQV6yL6cx5duvRkCaCh5T3YNGd9eSC24wFa9JEATv9
vCTODdYcqYygGZWXMdKlHHGNkMfK0SXI0uBxitNeZKT0Kc1qpL+DNTgrvsjUpztv
C+7adsuYb12kWs59CURaBbk+WVGDBqY7VSpC73KELLs8/szPk3AlqXooFfsNX8HN
Y2PjXFlBS5fgaaq8/KJhVkhDLOXsR1pcruq26QHsNI1hHf7+RsRpiso0gQsufDGL
tUPG55WirAjqmHUM4Z++s/7VJs09LFvd4C05gFDLX0dP5tTXbTKfQH218/cbJgti
ufQ/yRqaeWU3TKp0DbDqZaqL3k4c4DF8BNNznY2a28Hc0db8X4tc/tZG3bnImLfL
sYz4KTu0zjQjFXi0NYRNnk6Z4WOA3bekROLxzSq5ihHexFjQkbue0FoHdOKMCQmJ
kUbOQgsMge1JvDrC57L8LhJPQniLASAYB5jLVMlqK/JcrFF10lFU2hfZouf48Q0q
HaT5eza6SH+vAmuH17O9l3Eq76YTagfyfh8A2qFu7TGixyEu2LWLyM4zhKys1N5T
tbviiG/fWrN09kq+ChZkvagIKBMwU8G7vGk0dV/+WdjwRuy1WK3zsTe4BL41mc6s
41Yn5GuVr4LT1jDmdaEjXCy+L4UOK0XtjgOtz6KMLBx06wc6Zb7REjHD44iUugDB
TXCGaABxoyH6QRmC+wjIt+wUGV03rIyxkNfJsjQWU6X44tRkQIs2tOw0IlHx8lz/
Gw8VbCGS3vp/g+McHW8dOtqW2qwHGLH5CsIvrUKef5Z9M1S2YK9jAlDpYSbuwhZc
ktd82LinLuXM2KK/tMXiYmIHQpFSctLR5ky/CyenZD5NgxQbMO3+fUmhT4yZzpB3
SDCpp7wjPdMNEYniFtPS9YFyXFmzE6BLyB8leTIETUPiHVW4NRIrGo4RxKqipD8I
Im9MLQG2q5l5iaXY/8vUbC62CrshGDz67VAbBseVkzJ8G4NHep9KFYhuGpLprIT2
M3sPnDGtjWBTysayVZCoEF5Vsh/k7Asb+sAyFLi04xf5mhiiFRM64jnHFpboopDL
vl+NdiHVUrkMblSZUhxVu9kJoGp1w8GtDQLrf4tj3rOfGqjjHdt+30VxA7wNtrW+
GSNJDEB8fOZRXNdZ8ANVPJL/e6E3cChwesmfsRoEr6259mfANolIhXAC7fmhuD7D
eCQviBb0HTPrWUJPh2q9Kq9eh+J/KL9SE6IKdY1JIdPZjpqP8EM/N8Ky+LXcQcCI
ZrPERTBdfYLuSVa3I7oIcPvjzLJR7xESZAPJQeHH2Uhof9HNC0YnFcMa6M43em5P
htSRqBcbfRuFwXRPnAckchExrpuolIITha6qpCE7Hg1ycocFfWFnH4wT1hYPNttw
XkKoArT5YuF6vKrdTnoL/P9WH0Gagv9mxxMIarjLzMyGi4mr+o/k9sdouCW5QTH4
dekZq0vtkL0Akgd669u03AHTC958fKCAwV6dMWEFotub8kJ9TOY+tFk9yFxe+IMw
Xaj8x25hkmxcMmCmNQb9rnhozswfj/vkj5TaBeRkMfQ2QfA2Rsya1nPR1MQSqmgC
0IZn5B3j9o2XYzaJ/GkIHooqjcKSOv7XpizGemUkEVrdhyt2uaxSZbfQSdzTzk1E
3mKsCfd1lazPqxYE3e8TUAolKEsZ3ychxAxcgigUrJpD+GRDiLJOqUBcTq7hWiMg
07aZoJtsI0jeGKq1mJlBXCpTyjb/+tjUUMObaJ8qy5hZZeKSlHRjV/bYUjPpE1OD
5ki3cf1iBVFi/rm/uJiS3tTv9v9oeD1E0wtEZM5CEGIIztCTH9wru+vKGOlVXhd0
Xrw5qZUe5UmGTZmru0HzxFt99lAUbMiYcMQX4XwUxURDr/t/rqd4Q8HwMvQ2Q+uO
d/hE1XZr7kXN564PYV4jFCotLE8rIOoe7H+xxNNMhrC3oBJA0b5HMD4Fasbr2cDb
YWYGf1fIXYKQdXwOjHp/2ECMABYbkrYTFg66DY+mmHgNyiLo7hMgZ/DOaSW+OT50
LhD63CvcqQtlJf2NLiGFE++YWqE88+7x7dMypFIXrzcdkM8g5PPAC4IMjP2f1kql
6QnzzmejcN31lp6d32M0sU1yXrCpGliC1ENY2l9U4XpXZ9kQWi0JUCZOds78bXIN
A5bWCR6SPD1qDba++F0xrKVX8L7XdhHd3KXBUaHAj7hFhjsk/Mf6mQtPy3V/+hqk
MC8G83vUdsk2+mCTzXtQyXmUH2OJ1vG/99dQ3SY2JRkIWwEynvx0qnwYRtHXe4CG
TCwNMAwOZAk2Yi26bfnvY5/bheiuxe8Ee9a2arSii3WLPLhYaCSPH/b3lf5eVpll
UPmUF6WihE9Amf8C8lVFLCm1nNjrKOJANn3LgVo4OJAO+hB10rDP23jKivCTO+u5
/jvk4X0ie+SONzl0xTLqha9E0gA0k8r4x0l/jjJWHY4lyxcRW3kSMaO3GPhNaEe/
JY5BqIAGI1lwJ0G9Ln1BZT4ti0QJSw6kxBr4Nw6tkZKrwrOajF9GnJSgNzqgz1xR
3Jo1+4LLj0FrzCVN462PXpJOcApTQu1BR+lAwfNXvgA6pwVzLsWhVlc2T6fwNTa1
6kxmL/bzyseHpL0wjgO3hCVqFBEIiFb6zkPynTW3WH0wYgbcTneJf8JnrB+zu/zd
XmRXSjh1ei9pzGiyW+ZmHCbdVWuQZI45FwnADMZ0/XyZPxBRwbXYmB+c1657iI8p
8Z7HOMhnF3/EMMgXg18Ur3PeDTJ7fR8SWt+D/rqmdFwIsRuiPz2Wq5U9HRgJp2Xp
NAyVEESUffpLS2nCNANzgLcEuhbzRfAfFnNHo/05IRnxIbBBtpSf4wM4G2w3FNg9
1dLTriiL7VfsJM15XsWJv/AHye+tdkjQS9CbDekuxXDXleoBBVRcHCYMZsnmbyYK
dmesHqMzCcc8kZBqfEF3AMTDAUwZdpDN/b1BYYm4dMwxyhnDCvA1xvvGSyj2WH1F
k4xxdPHPIJ/q59J9LW8F3dY7PZ1tGqPV+/0Jf+AdQ7cM+wx6+fwtG999C4YEHdh4
frmHL6PR0n7QyjNSdBELAYSm8XdlcS/tQ9tbwRQSUH2VzW/AqRqGt3nhev65bNyn
ftBGvOeMetKssCDjiZv2frMIz42RTQ6Ji1WIcVtcY9+B1Age54XT2qeJsNX4K7vz
fUyWhyweMQWSM6WS8fkkDISXLuVa3e7b9LSi8jMCPGYNZvnmXU4PLRR1KWuyyrct
EE74jiN8gKpcFCkNwuQ/RkaPqnCqKCZjfEpCJ7bUPdsVaIJXrMcLWF0MGM30p125
jKk9IYIF2awutDIYwvWPM8gvbEQo0pjHyPCpY+2VAwP2PmcJu1DlgutP1K2MPIeL
xWmqLRkTkVU6FjntOmVtjDuz6ZRKKUs9UIXUMLVqvic/UcJYGakB86sgkCaGIsVA
7ckVj/e/i3xKSc0aktKOXXcxiS4yVCkimyVM7ohshjaxOuqwi9KG1K19k8VnmGY0
iRY3/YFvE8unng7k5eBcXxPicUjV3ZV+YQmTBzXUvVbDc2eBdINesclukvu/WoLI
xs4D8gOHWOvyJ4CqXbUg9Tq7FAkCMm6KeoDFJ6sp4B3vBPiymGjSEeUdv5JmX6Wz
Gm3ekoQYLznC+3r25GibkMlA2+ey1NecQKWuZLwN13gKH8pmCPwXTN1iDcFgbqFp
0uZRdyaR12dHAmOy0hZzWXAFTAEOJ0rFF/CMffK9aANy+xq1Ja/+RI3KtwcXanPj
n1i2IuGuOD0gYk/J/spEB81jJ9v/xNpwSLKGzzoj2erkQP7KL/k8eySyUM4vWzAj
10w+H3XQXoGGN5rTzcqhL4OBREZw6c1RZVLFyVRk0ircLzqruPy7KILBQCIau3CG
GCoVJDoEtEO4lhjD9AYMZU03IJq4KtkeWTjyANHduK0ADQrkrJtGVf580ypdaGU6
tfatmW/JOut8UnKgpjSCPWygo0PKNpNbAzAIES82EQ/QCLgCA3apfuxxAh5Tog1/
A377J0LFysNQts4YtRIj9F7U5CDPRdvUZi4Oz+ZbCnl4YcvWcSpn/0if1R6Ss84E
rwcMp6NzadzUQEDbH6nZ0O8X2lufg18r5I6ZKgE4W4Q+Qd0ASbvMm9vlMiPLt2s+
bTvh1iHdphSNw75kWnDJjnD4fsQNdMkUqQl191GylRUBrsbnXYcwhNDurK/BGBbi
2AVsBSD6AHpPZliur0slDiieEplc2IfuzZB/p4GuNYrbLHAk45mQMWNLnORYXlzG
2lWbveJq+kO/ALgLL/gyg35VwpYIonUaDHyD6UcJLO4BJ34cpQD4P61cJlarx1Uq
R2XngHyLOLZs76/Fc2U1wh5WwjzYqQOMBRmR4E5oaugiJ6SDs0Wc3bbxAu/tQYCB
X8XcuvUdbTqJzp4mX1EsEcN1t0RsTo2BImmKQmU4qdQ1mO/GoPUFi4dnTGi9jkRi
jeLLhICknd5gDou0S1+46TuwsRVwCLq9PPKoSg9X/crBwAp/ekEOoeLikP8wpCfn
ZFfMOPMi1bZbykAp5tKD37rKywPR4K1sIDj9gti+BA6g9TUR9hc0YiWxS/fpYbsM
mcbxvhMuytkgB399DGcs10vgzCoItS3waOWsIDh1/tcoTINXb4U76mzssi190epP
2CZ8wBOX+CVVKwe7xFeZ1yVExdGSg1cw8Kew5xLcmTBOvHYrpk4D4lS7A8D5SaZ7
uVM/WnHOu0OwRaV4JjiUesBV0YXsWE+COGAS8jjiKoFb7Si3UhSGWm0nWxySnWQ3
1xZAliJJhNVWL8e8rwgINRsSdCFGeVsTpyA2xyPsmFBvr+QfbwZnyiGhe/hA1vm1
sVtIXgTJYnmSilIyqCYCcXuJBg1FRBrUa2CfiZO1ZSPLOU/vF865O7ZFV4QMZuCp
2Lx3QnjC1dZ+Y7jFxMOdbrK1geKnDFgcPIMr+WWpSMZh25VI2gwyGvUbLiEa2bxr
eY4bet4S7Dz9ih2rZZQ+psovh7x885U844XCJj60ic0zVj+Iu3J6fqgkY8YYqD+0
W12VhjLc/HRzanydk9nbgMXSZ2MTRqDXg3bvpoJWDKjpPpqSKbFLbS0ntEEsZVKV
xJ2bsJVTYFMGL2OdedfpNo2Oz+IB28TK1D3E66VDoHqlGRDKrsWByKbzeeqmpdF7
/2D5VQ5R0GKzibEv7pBk/pAt61kz7yX1OP9yuHlj5unMxMAjtbMBODmKxkAutRh4
AtV96D9wrYRwPlktZ3qTbyVUnGhxqXgvEo9QIUygqhgiv+z82sWiv/O+/0IzFOl5
S+BuArt7P31Bo6J8hXXIwl/jojotFhf+I5GSUMluMxPs6uWMdne0ElvqIQJZaWwm
TeNZGLrCC/yU2o3GM31/1pyaWQvmMIJTILdS1a17yN3wtLqUPeOiLybclcOdFGFe
038CjgIHBTFQhxgkySg/ELDHS+0YDIMA6pJTLq9KtmG7Wsbo3CJLNN7wCKCCm44R
zzMpEAsPMMYgkky4dYzHC2PiyYv9b5lgyLZeb/myUfXHWdvyz2plBqeWUm4fuvYy
4oZRMXU2cv5bbJw5YJkplVhUjGwNFWl0ol5Ps7+xTLePNj0S0qnHgJL3w6KZ06ul
aLpAR2fv2GTtwoySnT33koksM5Lqy/XwsILAT6qR2sGofiBQZ40Ld2wpC+lwGrEU
VsfqHtZ57dtz9KidVlIYImfX8tW7oX8O3RPb19fqgutI0RKeq4NUxq7Ih6nYBrH7
O6VLzDkA6iFeVuvX5tAJEl6XfEoFsE0Aa2zVcmeNgWwz7UnxFrrFowKkk7oZ3D8A
a+piM4uE8NA5wIMpuG9L9n1OlNbbntPHEbgC66rnP9uQm14qhiX27BZ0ZVpkluXM
FfT8DARIPksRK6ADZ8Na/GMKRj3iA30HkXSJVQTg7VONrPK9DfSqTGdYp7tH5P5R
eZMdQo1Rs+goe8oEJrPtXUWgsw6xv8erdemqYXo7SEI++buRDIjn9pLPFEhHVuUt
6fOdUfgUPXRecfFAplEPLpcwoYpK3fC0VBMyIDxN5Sgoh8FaCGi+hqIgSDbSojvy
Spa6Ew4hXUIAz3JpDGHytOIp5B5HTlPA6widFqPvQoceI42tJh296g85iLrr1CB5
R9PpUtNtmeWWkTMxFD3WC7os+urGemX2VJghqBpX5HBr8v6HgQm08ST46cWOwFPz
5ODzHS8k2MbTVRambGUp3pIaOermvPKeGcHrbPnNesnP0P/7u3GfPsAo03WL19ts
Gzyxnp08ovQVYX1j7vYEu6usBlIbULbGtwgdGpT5OTRCdN5l/SkDRDnZL078Pq/1
lVJySDAmimvwIkdcHbzwb3GlRrwUofhDu7/Yd2zepTzS39j9EF9f/8wY5EKqtupE
+SN+LVwuZ7Bmo5TctqM640I3UyH7MaCtIYb/Tk3q3zPrSw/PpxM9TgTfM9B4snKu
BHsRs9MTFFzgLp9i1d5gcfVLRTaPkFvOZHYdlyL6DXRdJOGSNwIY9CvXG1J1uWkW
ssePp5trRUK+63o9BwZFZ7d8l47Se2YsmgDPVsaXIRYga+PJ35RQNJDPjOJ0ixmG
RnTnRHsHLMgmkQh0b4Zn/q9X0JP+0yhjDTPEHXU1DNzRec06OqzdTV88dc0PVBlE
BlaItCQC+ysIh7xKrD5LKwQBYWn7CzoMOMaENsbKS2E7Ik47ucQXrH/suNjE4FR3
VytjGYu5Q55MYzM4OP2oU2zXCjKI2Ap/Z6QnO2v5+MaLDnQs+pSzwwUGEZ8KsZU8
ZGpBncgF+BA+ph83z3iZmkXsO7718J4Z3ZX7g0YeJNIRu99sU9FkbXg2n33jC5XB
pU5wLnIbgunf7qhp/NJrX4Dp9OMwkJqc/Y7pX3yKxq+6n9hObCiKvai7hGhNVfb9
Td5n1EW9iYGeUETUs3ImpNdyiFPDYIpfFmWqdWDSsd6RGhkcDTK3owkNV7QXtWQ8
vXgQ2nATkxRytJ66cTGHMfM7FZvVIARHrwlZcY8Nlt21fPHbNFAb08TesdSkidrD
K9cf2+TVYPwRRAaGCTj/rgHn2bPzyPjUQeCsQ1VMebTAznYdjFi08s9T2HzLwfTL
lmVX7qVvPgJpy8/oW+/7sUTrmHlLuaHMra7w5MOOQF5iImuEBbMjEge1Z32UC9ts
vYWzcT/2tb1rAxfyRoMcrx2azIZg+s9TLlY5PJAyZpjK1mGgEgkku5UrYCqV/GEo
q8KVP/oOUpaEaGl14H245QCout3wzXqZhMo6xcWJaei39Vux6lnfvNp6BBV6hhM0
/BBYuu2GS0zqoUZvKLUxz6NcyjF3eH7S91/blda9sDCd/9bk8gO+oSudwI01vb1F
wzTDU69A5x9Rc1LTXwEXw1Jx+KvfstyCS4rzc76fpRzi8szhOu6u4PrE3Ak4WmPR
ao/ybJ3eHvFR+/dheUEWn0k+JYtXaucoVQ/34X8vHjmAjF2d7M9JErjWah6Ilzli
u6aikdMXojjPlGD9WVXnzviN5ZCVGio4wqa6mblrrgGlMXIG+seVT7BkWiob5/qb
4ActyQIecYcIxLjhhsm5mMfoJ/Aa7himXnZGahX8tNZGmGb5Jviaw5N0IeW5c0xP
oB4bCK4K9UYTmCb4538Dl/NxA58zSQzM9XMo4W7MaPZjEkdgrs6qPLmF989n/srh
4E/kQp9c26p8M/zTjhyoXgFZqEz6OxX9BgHssz9eH76VcGglrQcXH+mhehQgtdEV
sRKtUHdsZ3s+iHRDni6YdRXIVSkPnUGd5oHeK7YyyKRSDouuXd8ZAlGHgo5lHlWu
8JMmA5GNbgy7Oy6IsV9Lxa0v/2AX1v7UYgAYReyymuWYwdQsM89BA/sxgNFhrHnO
tfvaEZjlYwHQQ5hWkr/oImht58pmOcQVpJN4AW6nkSXAdnV7iFu0Y2Rmji3l2hrB
MYHmt72FHAebDuXG8cpGM5WTUaRO6wvIWrIBqQRooK+/WtZ5rLT3cVXza/hSqz/S
BAtsEPtj4g0Px+pcUPnJbXm1Xb1HF4rnvkquYcM503C0jEmGngl7eN91h1HMrhyX
EqjzWqqY7Zio9W0dwi1rHRg4ZoF31HlvlHAUUQzaTWS7eFERE0BXML1HPQVT93sV
3oLSNpYb+k6Kvu7enMOtELbLWsQ2FL2GogZuGTH/1yYFJBzsLMCJnK/y15VrGpuZ
u+N3c8MqTb7d4HRVnauwpZOh8Q4uN0Fgoqh+o4LifWzMFLRTmVJxALbRMJIfmWgJ
Qb/51JHGg+E7GNxFDP1H9h9h5v/+OArpqamDMnkvwF0bk+FCMQfn8xFRuWREl1tf
mo4G8z0S1HXCCBsrMJKo0muIEJkfYZcqUBnQxpNMeKNo2BJIMY5hJLA7kxQNLRfm
Lx/wIft9XwUyQaJe4ZrGDPtPRW0KTFfr6NVoACs5Y7iRH0j01nD50R0tF50euJH+
+391QYEPpRafEX0B9m4oyTYo5TQrMd2PVhipDNRcW3oslg524XLnwArt1EjdpgL2
xGS4AtxD9aH3dRlaxI9lqsp0lqCkXOy24jWEpLJzJfUqyOALATFv2QDKo9W6XNq7
Zs6zRm8V6lECfVvAPZ01wCXRVErW+cGcnxDca6FqKG6Pn4DWvWA+kB56d8XoN7L9
GWuRFNSLzoDxs953nm4d+sstA/HWlTQ+n4MRHAunGhcjByNo3YQvtsMc2Rm23shx
U4v8DIp1/6egirQAGY9+HYyF3BYs/9P4dypoUEl96K6IvhvprGd4Xv6zPURnKhhW
8n5d+Di8Sg0BBG66fq1MUtTiHjE9geOf+OOgNoWd4KxYXPMOz0o72Y9ZnVExm6QK
e8H0unhilzesOLdlcKwC3YpLtLuNHVpfu9tWCh6TFZuH1TglwBiudw80a7yL26uT
KuUbM33FrEkgGHLAlLFBpts028KggMDAxjdzUkgAZryjuC2KbN6sQ9RWAU9WG3Eu
9qrLfJaVwetMaEtGYfCS0c8RfYSIqO7uEUsqPHwQ3M8z6ItLop9zsRu4YM6rOU9y
kGTTHN+dQeBiAo6VNj+43ia0H0lXqukX571Nq5x1/YhcAX8Rkq/BChContGNFCr3
AJ/lIqcslp1plKAWVYktK/15BBYFJ8rXtgN35mb4/JZTafgRd11xjpYtru4rgHmD
T50nxFMzO7hmJCyXCROHZMqxqa9O0p1PHpJr84LjpTEhCks6FGod3j7jnrDa/NMo
eKUcRQ/5BnH9gLr4cbNxkWyl7BqIz6mX0zG3x4WPtKKj0tEvD9SOoej621LG+IQk
mjTJuqp+YZG6HbQXYtbQ+ZCAnfTjsVgVdWUN49S1yn/4FoT+tQDNSu/X0gD/jlnT
xQbQmHC8nQ1a9be66W+Qapbh176eIkZaIV51n+Mqh/9mUBzWUGBTvGQM1d72qt+8
cjpdxmMFsBkqWmbkE9dvUQLltDCmZnuX7zLilfevTcgZ0bn3v3mAti0uLdM5RMrj
ULKWKDvdmZ/WNkcARYU8Eu+kKsQrEmZm6O37HNP27SKYDhUlspuCRKf+qnBFyHyv
AjNsQ79ds1Fl8/+bEVrlhw1xVx+G71sR99rp0m1gdgV4RzBw3Dq/ZGvBvsHO/WI7
jiL8m6AiKewYIcM3VUg+eDcAKZwInBAcRCrSSiobZDZJr9df92jIsE2NA7NRZYqa
dvJjPuqKvKNzxbpm5MpgAjqj9n0ePuPpfnxGdFt3UnXAkDaSKE50foIeG6jApYXl
lW7OolU0FkGBqxNdp7moLSjNmcYirXnTdrsoIBkG16uaqnLEoGvnIR3Qvqiy7dW2
/nYGqr7sdYpFse5gRCAZaFTC57jUuW24ZNHrM680sKG362k+QsORSDzQljMy29U6
x5GlCI/IGtPqw/Kt9dkosghDOEsGEUJZc6AKu/tHBBd+NfABJEWazAJ4TI985rnz
0ttIUxlScyYh4V03uDOY6nStSpgsUpEbW8j1xzmJ+bps8m7HMncxO6z4YVu+ZWPe
DZ+OVEMI+KQZab8v2tYdzDmkIdvP1cms1dQXi4Ow8xgvfFDSMnzbQkuddLrSMVkF
9bqOpb9IRvI6Zmtte/xHAzagKXdJuT1n2TSXzLWnLW/fF8d8IEEAZISSjc+i+Rfw
7agi3jbyZUcDwWSYecEDVnY4BiM7l5o4236OkSnsuk3HLsKWUZxM9uxs3cylFOJ6
gyYZ7DMpf4bawAfPNgCkzvgEzE7xkgge+cpAl45tA9MhDI8NvQqOVbINtdEb4or1
uyk+jW3658g/BiKNME5R48fglO0T4lXtHRyNF4J8JOROXKbfqxB1yMSy05TsnjNF
8dJ5RZtNPbp+xw0be2cj2WIw2c614lSK4Xia6pbibr/RpG30AtgDsT6H/tGPmWev
tr6lCR0HeVhPsD85I+jtXFOMTJV/JXHue8NJUFD2nIEBe0KbMdGSV3wVIQMLFN75
sqOBJgvq5qn+0zkA2yI2ztJZtTmxRNKy7PDuVoxQimMB/zH6WaZcPvrcyGuvCKga
ejfYzN+p39JmWE3sQ9DN8XJwxv+Qj26iLWBP84qta3VO0w13k9EplRnS59Ao4Zwn
Xo5qQ32Xqx4U3TUf1Yb18KqGCojr4IuhVn/CEj7LTRIcPTwHHJJunEmpAeTQmJgy
NH17g26W6U9Z4zVO3Xqn1QPoCFnTcgylIdzSSSfOMixm8fkfBlAJVXwl2df8aTJ4
cX1MoRIf71tQ2lqJGlVxpP9mSLQf0dVske8istw5FtrdADEbjtlBcHNqrhvx/XUT
NaKTsTgDoLbgQWl+AAUAH3lrCsh8v3fQVzubqzfBBBrY2z3LVIcG7MilahCm6FF8
YBL+vaRpuewESQmqO64u992c7KBHS28ghfvz+vm0xSl12BjNv9aoMxTLro+j3+Gc
kF18JcObkWiAbdE/pwl49FtXLAAkxQ9djppZi6ZQDM0u9eKKAMzz73r7xd7PqkCX
tk62J68dt089M9A9R57hCdU57+7q8jOy1qTU/eD5wYR/vsZkR7c472gUsCA93gmh
g6Sf6OMD6r/pXFxQoy/541GBjEcveA0o5zCECcui6HHrkJhE0L4FrGV/cpVQzVRG
Vtw0KvUq7YQhNV4Mkg82SOJCTQju/eTvGYl6K67MlfvtGE93At7detpNq5XjX0sj
rSDLFMcxpiOhmiAIEfI/PjcmoZDwIQvHZKfuDxmrXE8uSJM076V8bmnwGPuMZr83
DBp6+5MZ6VjUyZyixZb1jOZqVrn0mmOaNJjt1+5iwd736NAUmE071rfP9/PPpez7
jiL9wtJUg00oV8BX0Gw5n643LmhWpcdQOQ3GBY3ZpuZwiBlWRmZJ/PAHrlQpqGF3
B9/lmOCQD9DzZ8rFvx2PPyLMgNCVVXscpRLnmSLSlMG3tdFw2Z4sC1zF9RQ4nPud
xxWqbXXOLWI5d/FpOE1PxCKaSRggWkHOqq2ama0HS6CsqCaeQl7dfKyxxUdujnLQ
frTm1d8jqmRCAo3qWigzxqVJaPCvkCSZOp5UtVCXBPkseAAYFEI6OLoneREGgbD6
qLACIcgVzFCN7aYIwcJry9XGVK7mxwl9zgGyBAFRC1R2yB4IP0sX2Fu46Kc3cyX9
vVHK5kqnUV7F/UXLxY+2qGjLmYFsMvQGZqcF84650Wh8yYtLOB9ZlrqFatTvcc3O
kytGehSqT+rxtFLfgyy1jQ9wV8hSLKjfIBFUyvLtlO/ELMsXyR4biqd3BLEZ6Tp/
ZdX/8O9izaRKTeQn1HJp3joufrkY4NPvc9IMu1wYWs0pu4WcGXvyRciG6d+EYee1
39DhjZJSPBZYGoXNk9kZVJXdKFpR3SOuivRM/pgW3MbBqT0Y76xNh1R6AqdjlfbZ
eGL/fmr6+TxEU61mSBdWOyw9y5HPzg/YzVZLD0gjq5SeGI+7OUU36LkydJQZSpqI
3MhTnlv5g+Nj/3aUBfeUrL2M1oqDHSt5VfYS+d5y+R88BJ1bewiic1OISR8kwHMX
1va8WQ6ddONGnjFmGZNrWKJTjxoFS1JXb3Hi2ylWMbIi9e09DeCgs7LRu2/jEkW4
LSaE1a5DD6QnKnyEKZEfd5EDVQk7fWew5TEJwkqCCHb93dij03bDqcyAQPq/oV7c
eQXVZJvie3XH3jKABB+oA4mK8nl14fPVG2Oz2moXSGTVNQrM2HXYHREMsy6EoriL
Isrvm++UiderD6m4V9N3/UokOoxMMejpBXV7UCxGfIrUoSUnHICv/CvJir1mjWFY
0esPHMNWvRctGpkNR3apEF1yAepeQtsNcpjyw7i+0fgghzf6nO6KMmYi5skPjdQy
aNRhBcLuyJ1pqj786PWY9MsfazqYd+zrLMXniUErpZNgeeiXzsvE0W8XWpn80dWq
zwbyDQl8fvKC1yzwcm4nSeXI6g8U8TvJDeJ1v0BflNHaFyX/JSovNhuDxLpwA4sy
74gb8fLGJ30ZmCjlSboaOoAFEo+y/YUNqcOoPKOBNPZKuIv9Xgld7sm8VgQXZrjW
StIhB0uOPFx3Z6nA3uTSYdmXvx/c6lzKjhvCdivZY+VX6DFGd1VH4k+Afez93UDo
97q/oL2H2uYW8vNastz5SzdUG29aaIDmdK95tIfvCrDn+IvoPJgSzdy4A7Z653rX
6eFgSqnCF2I09WIjAmrv3h4REGQoud05WlK7VegwbT61vxiqMd8XAPEuMVjmSsBi
QnOy/Ee1Op7OURo/4VUE3OrS79R0rRFjlTE0hl7mowh1MomLa9u/Q7BZZipsUFGe
dM2lZiw4KAKUMxzsz56tXJzRZn7UST+znotxzZG+AYKBS8t3mSYdjzWwqZ4yowCC
XBBXO59DJObTUW8eLZde41160cWR1FeBt53RKQVRHdi0lkuB3KMlnEZ2zSgT/K1I
c/u81nGDCFkA1SEeNMQiQrS+uxNZuT1JbPVbmPwtGF3BDb+Th/nwmooRMBFukWC5
78R35svyrkPdqbA0WVhzQIZNRyz5qunqtML8/tEa4IP+pXIeXLQzCDkiT0IU0c+Z
IgCFm2iOuScxLc+QTDhk0S7QzaMy6Y5PiQt/4VLBKA2dxGO8Uo6ptPKzs8ZqF/hn
Y+C2ADhA0fV1MMa7kgN6gUpxkmKv07jZYQsMJCY7cFu8sIgOuf5TdEgQhSgIsB0I
UP8I+3GTb2ecK7WWYOFV1LUjmuObdfn60kKuUZbZ4WvL3GtTZia/94tauQknrjcf
TZ5MHNcCrSe7f03dcLSECbE6sHzR172e/5jW+PhqIzN/akU2bhXKDgCgs2fdBLFA
aSUWYAjJu1LyQnowARo401wfdM9N/TIZo5AW2AYykMZJkt8SKNXQ6TWOxvN++9VG
u6/g7ELavPidfM+/CJ0DTLYHSt+Z3zKoG0ze1nhtdDHLb8Mh+cs1aWWiEW+m/epg
RkIKK1ybmp6swduHLe+gehRSP/dEI7NGUMnhgkfnIpqjFbUevDQKABwH86hugRth
BllnpQozA3vKgJVa7mNmztmE3oShkpi5seBLRVJTaJkB84Fim7CFuHrQtkbglmnJ
eDWAabtRG5dUva1wi+Rm3Hy8GfkTWbmB48aE4gm2q5i1C5c53Yirh45BVv/usIAM
WP/LgD2CAEsLHyFBQaRG2LqTs9JR+16/XGhMtdb4QCON3g0GDoewHHo6P59HVzIP
WPrDcgEhcL81n7Q8vTMxfD8pmuVzUjfi5DYtN/8pTthxWRRTgw8mXPX4x0Qq3tKF
IebWTKrmveo9YyKVjnfvR85GWHkTxjrThufCu036T7uio8UY+mTVm6yiM59LOBsk
hU/oT3Ue0Cy08EtcQei+2XvtVyNis89LT0J72JXP163wEPyF0C5FLZHOkc5dn8y6
e0/SBF0iXR4IVdlJpSwErIR4UJZihEJb1nmOnFifRilW2qtLVptYrOYjHzPGFMOl
oXA/SsuE1+jddADmQbbOCDFMUrNdwkENWnpwB7YYViUTZic7AVif7VyTFCjEYuhF
NAz+If53ujUxhHuzvDBoKBCOoolSv0Z3M0sFFZkTaSDC0xHqzoItrWW7u9ClIW8T
IuT2vVAiQrDLjh6KMeLfQ0tnNYiHKQDfODIB/DHRiCilLaV9el2x0Z42Cce5BK6o
FNIIsPR5ptyLWXdF1WXtMt1/yJM3P1W9acreuYRmUoK/UmBr0vYC057QPz0Sxd+M
BJvu/p91ZNKhhK6JnsqK2ijG0Umt4+6JWlX7TWzB4WZfmGKK71syaWxp3ifNUbUW
/HHAXRigGr7Wu9mUdtK8PeujX3B4fNHpdUKX4h4A9ylaVj3YjFQE0EHqi8jwddKJ
ptqoHmbmVANlRUxeZgTQ/bd/thI/iy9x1kch2eIW6GE8x1M3X2T3yqZCbE51Dcpo
23nxgujxJmHprpBQ6nnqc5MSkVLMpU88aBPo86rjuVHRjtFSdY5O8NbDc/CjrO+J
rsKHMKroiOV8rwmAxLtTYu+XkpM7bHY+mvFYhVTKIHaQ4Rr/BZ2YrWkgb7l5bcA+
8jzozkx/1ZnFxvk6vzS/jE6U69629yY2p7UFii84MiNuMxqwcIthVJxaheWoPvlH
ZXw4GnPHR1iZUZJu81FIACRIO8RH8IT6bsBXtpc77HZL0rvxFUUJ/YVl1MEuPb0f
VQSsJqrIvK7ew5QpGccLakL02HdHHzt5+hH6eRHVMpR1ymiImNtbCWBTpC72bmoV
hCTOfUblZQ9meDU46FjIFk8JlgcD2vpgRsOJDREKKagLdb6cKrqPWVqKFpLaee7s
XF3l12s7Zw0DMLpi/7nFZWVfe/KO0RtJhgttTuuEi8iDwzqA/9O25sNvqrLt0ty9
KtQbxaBP+mlGVeFXgCTVkBCDYTLLp2rSmKztdd36udGGs2Ccm9KTuvsOAXBmSykG
VDLtiBhkxRA66rCDSg8Yw0PtVqpRsrUlhc/ITZLKhwZdSM9Js9x3MePxuJ8gM608
sSb1oGyM+4vdBKHeEE/m8ojt9ft8ObNJewAUCXkgr+LbTAa4ozIYlu6Z6vsklUPe
eWZ9mxrt8bvBZqjKr93LAOMWYdTc85ll9Gmp/FOFg4k3xB1CpXcSkBFNcgeo8hQh
agi2NQR/OZI0cRv/kxf8V+NBzknGBtNoRuE2fRd5gol9cTNrLU77Dqv2J3M/Y8Sf
uXcbS35egekL2TSwQJWJzTjyXxhyo/Hh6W7TRwERuNKGkeHG12ZVHfuaL1QlzaWd
ZQ1aNp3eRH7nQzjvaWhzH+tyuhmBmjuwNk8sL1m9n70sHfROjkpRQoFigKPF9lkQ
NOG7ZJgj+S/gvJNIDNG6tTkMdGOIYin531yiPOS/3zOTiNGFpml5BdFQUVHTQCSo
DWC+fc7ZF2gVIvWCIlI2OEQ22OUal3SyVFoVED6aAfcMk5LlbagPjFH1X4A9E2AU
IdlejDIdOdyKTjdLZS6Q7TI+dtqnoPfRmd1fwXKKah9gwrRJVCQ2LLzDe/86HRdC
l8/Iobu05BAu5SqAn6WIfpmG9edpLNafAL+kaSsQCmNWgIMqp3tntMxqRZkT3U/r
X9jJulVqdAF1RvyukdA/4dLl7taH5JAjxKOLZZmJNAlAlHtlGyy/ZJwS9PnFR51O
hgMpUUmgNSNiNJ3IjeLquY4zNr8NmfMDjD9nfXm7P/7WN+yok6D2WI+aHe2yR/W+
J7fCJJRkCQGUexMjt8G3BV/lyF2MswkWdEbnH2Q+NrapuMDD1fA7zR9gOAS5S9qK
OT7QlilzesPUaSs0pf3Rn5OQrf+lwgKpBM05om8nzb+ipBsb83GwR4i85CxWcjZO
rF3YqcCCqk6MZWo/YUz7tfhBoDwlVxItbx27CMlF8IZol51/VZdvVbozS9F8iU/W
5Gc986/9rhUuoa0cSEEJum0Rr37el699HlKfjpfrvH29UhPoTWuac/eLjWZ12UnM
ywY/lKjBWpDfvEf1D2SyFjO350JRy1PDWSBjTzE7QUpzr3dlXkq5h18pEA6+o1FX
OpmLfly0/iINt01znRs3kCAz/8r9h/iQeFMA3oCyj8n52tiB6BiAcHzGebu9FQW0
A/3mTnF0aQh6KrWzWToQisY5cdwx4iHlKQ+ChzAsO2ODfRdxnDUkuQPFCNLfBn3G
ebT/6P3nOsItTrcsbhui6hiT36RytxLyUl13E86nhqynPfBsN7eALiHnGA8EqjNL
O6o9hvfghOpS4IN8Yo60GBq5LpZceqFK6j3LukONH5BjFxSPRoX3XUDcObzi2htE
2t81JOrKx9onV1uz9uaEAgNUmDu/1PclULd82yZAlD9vsvBcZkPS/CBk1db1mvCb
J3Vbrz+rMIz8UN79kBZz/u8vU7ziYt/1XOXVSc7WDJSefECh8Bwxz8VJ5liD/ZoG
Jw3aNwCEnbYpWo+p+MydstPFDUkTdcUxaaRM+UK6dO5BfCgH7W1lUnsrRwfOr9YO
duxEmVK+YqDWLjogdS7pKKUC9rSG3fz2PrNLo2SVoU1LA31zjZStYcZlLvWHWXp7
6ZP2STldYYLBpqirSz9kfwbtru0pZREoMOKjCOXQ72bG6TAIpZmzqoZyJa6ggNJb
shJtz5RySUdbtfD1LO/0gbOYN2hmiFEgodN+2je0A5X98F0erwchNaRdQ0Q7emWZ
wUh/0doPs8WHRWhUjOup5/BshYHZxuyhvxHyOCRMao0RVZzo3ZCuzIq0D/o8ij9X
MRED7p5Wepc9X8JiVP7ACx+g+iQ15I7zTK2SEiAiE/qc+IOUqcU3wcvq6+075XsE
vq4zvg1muelJ1zYDhi4A5QpJKXf514N9LCS5OnlVFGHFgqXfsnMnxFfvkOBrywfl
25Y5J+JeEXEo2r/05saVQPKR1lUiZ455tadFVP3pNo+wkTtXf991vYiUCq8Ao3px
aG41FSbp/WDHcKPqNw0MkXQH/D2Y/m3Og0VjCn6bZWLv6lucBNXKEG8KT1yX7KRw
ofou8VQaCVsoeW6qoORiuo03X0LLTfMpVK0q+/GAEdt/HwPcLV91kAatPIBGJC/O
rjqGz+pUW2NipjtC1q+YWTL6OZ/0HO/PkYEGaYn0545hhmRvNKRXNE/jxwR+wyB8
SOALvjUJJVdlagSU4XNyuDESjHf0aiO1WGYymobbeRRZFuAB6fEHHLhUUFqoc1rv
hiPZCEOfro6le/MfYrfP9f/SPZkutyqXZCVJ7D3UFd46KD6OZLzNBkzt1CO6/0bI
aF4pt3Oq5fdoQBVht2d34Nny4H5X1WHNrcBq6IBIwQsR85taBweYy+IIOhtmWdMF
xoCbKWHGob0QYq0j1AUvzmI+K15HmK3/a+4pcAPuZB3q4RfSpddGMJPgIR34xiNQ
GaAQj2M6Xb/swoQAAAeOpkahmdG8CEIaco5J8uTa97sNUe/rui0g88ShnjsctDc0
q5z/R//7tAHKmSjrJhcsQKKN/CPYvM8vmhcXrQAzLhPuBpDE8j8BnglhaUNAvMlZ
BjBB/JjTOEXgm+ExQz41+YxremoIa+DuEjeKGoQRR4cvTSAb/mR7N2x3wQQLwkuD
iM6cKl4XzSNIwyWW5y5T84cd+46/60n94rL491Wl8MdMrVZWUtgkf8GCKU+JHmhE
8+C6KVoLZxpmuWDBu22NOaFa73Q6V1K3HaIn0hniAdLvwwUbWhvOx4hbyqxkp4h7
YLyOcCNAyV1WQq0VvV9TxBppOy51xHadsSksEyO6A70wClzNvFIyxtMOE1+sLHuh
N9BmlP79QcsjRwOFO0vMdWjL5kra8xM5kE0H70gUGxPHpFY6hiNwluM6DrOMeHDH
zS4MPEMfiXgjNzU5suQa8TN86tlu7XACiZ7pkF5ISpVwSGftoXFuIZ8n0oM5TYM+
u983F006PpeW2EFe2U6wszvjXWvsw/13QxqvvwPerkYvN1difCCScJUcMrWwKn81
ndzDrMxmf51sCLAA5YQXySfhN+QsBl/FZ9JE8X6Ds+wRkVMqXm9JWInL0E6GM7UR
hBODJAtGWbUgq4wmqHoFhn/cR6Ykn8JX2gGbgdxfTxMFNdPsh2yqqydiC/Nhd2Lp
XyK2nDrPYT+NQ4j1gYrmZ+XrSlvUgYFBeY3XnBqnVLhhYjjowmiTkDOjhefNe3go
FioXSFvlzklfk+FuSlaiNZ29HUbtZzb9Cu2Wol+aIo5ZeEH8XEbgCoaumwzfvExD
pliHO6tuR6ulrdhNsU1XMgyOYoY/1+XZPwK0g4UPovhzGIhfpjbjObMZOPPoiTxQ
QmEwQYQ1w6G40sb+I3epEPiBw6m/6cJ+hHwZYFsY/nyAm9fkIvtB14ckkZROjKRJ
HoNZ9NCuey8oS8dlQItf8EAsfd9OcIICk2BDZK8PGHLdRxq6JVsxjqNWnPSrxVW3
O0htJRqNlRi6T9aO9qLSHEIx+wylSAOBmBwl/VSXHkik0CfzEqY1BoBfW7Q4OWpK
IHnAxOiGTx3timz2HRyAU6DkpgwK0PexDbh1Do9NmT8GUCLYfie3kiOMTm9eJB9G
itq5KKgjHtv4rhtAh8lUjAbGfigS0h6CkI6pOj1xRALIhqxBpeXlRp6q74V8q4ey
KuwJa/hkTpkTk0kt33K5crFaXbgq/cTZBUZZ7iRlWQjbLLIFAF/1zKCoxMYn26IO
xipu1X9pOqf2j3njWxgRF2/KACI3NRl0s8qqR60WkFocBdSKX2/o4oqiN96jsLez
PDrXqyo9WHVrSqylZT9getvZ/r+B2a05s7ikIVrK5EkGmeqU7w2qkiDoEVxhxwO0
qwh027w7Pr/ykz918fY3yu0Ko25b8Ze6A6BkBvSNU89J6A1RXKYSydkekKLhRjz5
6WMRoH+w0aSaXhxdeK9K/1xPnhJ8AFlGkW96VeKurYgvy2TQMk/TvoypfpdxWdaH
uCfbdCi3UylQF7FnzqoqM8jFSk3UL3LNK6qsL7iUcdfdISYTOFkwsRr0fnSep0i9
3R163LMOobtV0PDrJ7YVuRB0Pbh19djucSxm8mPSEySWMMblaGrMHkle+bl6ADFo
VlWxLBIenwripx9GHuv3YQp4TBQu58BjQ6mpHE52uzZbRDQkvxGwNiYtXECQ1rhy
zeJ7Ned7Y3npHD53zE1n3EPsDz3mc7OeNQ0DHrhrw8hSvoPEUgOQhb0uv5e9PP/m
0gDz9de87ZpwpeOY5ShUfgd8s9f+B8DCAVUoen4uReEYzkLkumP0OP/f4+yzvTqp
itxVpCmWUMpr5aMXMs+0ltbhFc4jgItXwjIOPoQYWSHHV2z1YJRt4pcppSe9dR8R
ekkRcOICuxZE6nA0lBxXJKKgKKV+L8ch6hTpv/iV/4U/4bK/+eMJ5m/Av3PAlGP+
44mwSLuw5b0bGH54jpuTgy7AtmMbWa8+P7GQpEfkqCRoJ7X5rSLTWKLY4rdSczLQ
PfHMvumnDO54fTEuFlqbKu8Aq4Yb05hlp982VbhfKi0owfHgLP038dtzunT+QOM1
kdihKlPVyiwSUhEAktF7XNX7QdB+p5Hn6oNtZsjmX6Ybor25Ja92RGXxcWgBX9LK
sRKrQQjmt8UbHf9xX4NI9/BzsfhraahlJDNvC4kBQQ63sCkG69FxYiDx1ZkR7J/o
o60ofPuX+ZVmCLMkiFI1H8pjxHN6iMBaFj+2TbAqnFFOgT3CvMiqlXomg/DYLKrP
efAtdn43GJAKOyb5btI4uQxkd+J/xFWGGdqnZryHQjA1ktyXwhfQLnloqVEbdZZS
q0lwem7PgGYB0nyH8DX5CaXiLDLWgOyVj1U46d2WPAq/nVlQbpH156JOAw1hvXd+
jbUOxFqpgqkJFgmiLelJ0riB0q4WjaM8SBRpzVVlSOSyZfPUHTLrV8axxE+lsQc3
u1fp0zv7bGmUz2hacihFhU5undz3Wv3xKqOa0LvfHj8c6gPVKpRl2iD7h+2aj+6+
md671t50p6FF4AeeA3fYvHpr4O3L11fphiNDyI2fbax71UD7PgTbAh2gBIArdBh1
m56zaBAmDB3ofjs9OEEH9M2YZHaTTEa/pQC0jF7jPIZsdxKqupNTR29VtCCuw2Xu
VHZFVcEbIXKlXTGIkmhkaqk5k494KZltQvWVd/By8nGPAK/u4LHpEfWd8n9K0C6G
PPrkay9WYRfIjU+bO0qjLl5Qfmrr9aAQdypKNiAogZzcjzSgkAENUWgzYYfI4eJT
C5O0W/DNzs4U3SI2LbQp8JD+S2xHT2Be5tG2mjNRYgOg5YjtlftE4JjQbyIhrRJC
REtdnD6lYHYE5bXCfCCztWWTOFPFMU3tHqPyA4oZYekvqAvG5cYFMFno+JARluAq
kzruII1Pz99JqZdj6v2ypidh4B0oRPOboEuOZoiB3i4sxTs8UhgGhegC8x0AbG1j
V/Dl73ffx71yuQj+23J+sXMOmGY4kIQi6jCo2eGODQnauxqh7cCtwOqIKy/M7BQh
m3KdDeQAryePz8/b+6RAyQ0jKosOTWiMRApLylXNj8uB3GXaRfTS3vd6mwFLw4Iv
V2xGVv5ZoV1p4lht5LjvTLP1nUkL7+sbDFr3yDb8ZmXQpzCHIZ2DH2QsiZpwAACX
WWcJI/5PKVmezco8EyvNuvs8LnnTKnRXrWbehLd5j0GqsqEKbj3kpFzK8Hb1cqNH
Dsh7KbWLCd3nHmoWXbuHOpUbeXSaejtIGu2Mt60sRv7YZUUK1xuyjjrvG1M1j47I
SQLLqw3MrpoQKQFnH5zUa2S3RnpqRVnWV0xnH3AQy1OTtKsP7P+FkYtilzkjflzG
88oFSLvX0oMYQPH3C28+dCXVsyDHuHvTkDFRCwfB+cTAAGHHflxymwClo7HnCzpN
BN7PN7QCuQQIJ+uHdo8QTtISWHXe9ciQWgKkNqwC/h4OJnMN20LHbYDlO7xBt5ZS
2XG09T4tcwF0/2vJKNu52xoJg9iUbsALhP9IKRbNZoZwAqklhnj18zpevCnb+6se
FfS3VXH25Wb5KXH53i/2jqZc84YMCRWWsKj7E3ubcjNTSoM8yDstzL1Aeb7UizLJ
YKEDqlxijZjc2diTFxSSgTUmj0cD9s/XmDCvP8F/mLy2rTb0fdoPXNCyQnTX+PP+
FLl1AFdgKuOhs/Zvjzrkukgf2fwOrt9EtLfse2WWYlaa4+ngu7w2TeTzAIx9LKSh
cO528/hUoXjNxxmbPWpH/qboCy9XZFTG4y4Aqoa7uyL/xkHwjusMOr9y7VXdbSNM
NKSzcnEPdgyXx6kTfl61szcOZEQGKnmvy8/AbqLOH2ZX6PfLR/w4PHWyH9ZE5EHL
OuehV9aZWEt/Kirw+Fsuf9VJeup94A/oYslDMugeeDvBiz22D4yFtQ4GuFfcT4Iq
2IVDsBUU03rpuLYL1jIu6YbfB7ClSSRCWBp76tB5ugudOKQ25qUpL/aEZ3/bn+9m
Xv46uLiXNOIUVoG62EORgJLT6JPyXf7TsFK6vACdCUpEq5npVS1NbaQSGKSeulUa
1rlLO1ivzEETiX+wsw0/1y4/b/+t8VkyL1X7PekRbdE00jiU6NSbld0fXs6KvQz6
M+16mmGlE4rFEa9HOaOFJuRL4wGr5/9isi9oDDXZRZ9Ogf972nsttrj87OM+1wNN
asVJYf+zrtcIY1ynaw6kK+XK722TVXINsEBmwzW0JnVsd5yXs+Mm7F/6AB4fBxXi
PdXxPG6+rlMYc0i6ZBNW714Nr9HYRXVrWyw/myvfo+8Mohy4qY11/znxyGGd24jb
4mAUrspdJykH/WJpFSFHRYd/2pLuq8ho6mf17KGHA0vP/CksXkUZ4QJSMUK0Z4xD
3qrpEfwBZLDXgRDsCKKEvpZrDGMKpJI8gIrTkhibhpJOOMhEHTi1KU32nS89NQ/Y
z3PSxdY4r2FmYSnSU2+YEMpKwSle7o1MxkYYsIOarbqkjDVJ4Acj1gSap/+7dvx7
1iPPPa4VfJF5H157EwV1ScKTMN6dDmIwQeMWv7S9dOFjCCpL6Eqlpi960zEJLeoc
RAF8+T6NGZmACBs1a/8BbpjfP1g6QQ1C1pNxfQRUJl6WgeB0PYcSNFmr/aYMj6AO
NZ93HmfOyHPipUQitfvjvbskwWfHrSPJK9FI4tXHsD8S2kdAFbc/MOyB7ayAKhrQ
w8KnjTFP78m4M9o4A3FqK6psgrf9LRKhxwsb1cuhzTSCkBGJ1QCGTIskLGl3sraT
TUMJ5zOMSBUjN9r+5hjo/iZdb77Bz+eVQbzJxLbWM1SCXrQDwlqx2gmCv8ZAEDvi
aaZPEbrihOEWNHrqnmw7wL/Xq6k01TbfH09p5Qbp6zBl9qzAGIgKIIcNT7Nkm1Dj
Xv5TbLIm3FmzYLFtDvK91+buT05M0SxQWNgxyFNDLlavsRP3uOSAwWwJT5qUJFDE
bY/iK0hfQY2iJFRfhU9XrW3cvdbQxRk8sPqJ4+HPFrDqWVa67Oiz5LPDlIC+FmNh
mJgPUZCbuv5my/+GdG4M1gEqH4Shyec4xKMyQ9TNtVEXymn98AQRQ0Thbg++fFhq
Fs6/L9zN/oX9MQDsQ5AQuAufxvOKPFwoJrAqNjPSpvSoBwt8yEmHq+d6++J5Qjtg
ysiKhEF8xq6v84tYp/YTZe8FJUvyxWbM3OAu3sLbYc+mNNSRv7Cfi9B/lqrNmBYR
TlfafnnlrN3W09tNaTpfK3akW2rKBPhKrOWJrAOad1K+W7G4aVdzcFZj8PAvEJ0I
GZY6hfoRete7a5v+ctUFkxbZANGxsbGbq7sY9uXb4NHlLo+srkZp7vBKO5rk3Awb
4p/tl+5c1s0TtcfI675zyFDJUFySbYmLo/GJ73Es8c2FWdavuMRfvxfvYIazCe/B
HyVEOg397t1BEbQiPAErZotP/5VRJ+H4vr+Rb4rQe5KRvOqkEhG70eYQOX9J2fBz
0R52pQfbOl9bRscdtHkLPtUh0EhAUcydsg9rSJW9EvNNpN8swk3v8+xS5PJ3yVMk
1UDhetO/G+j0kCXRwslz5vYy91vah7qQlKims+XI8VrV5UOgPt5WyMRHG/kSm6/j
BuZinniqiGhDgvCiku2woley01q6JvCPlaiuUE0TmmT+/7cYQdopF9qTM3wp2o3c
WGrOGIhJOyXvHoXEMMiWFIhZl2Yq4lRJPr1Xa8Ja7GIH/XEhMLJWQY2NoDfl9mFl
zGRT0WSNrwu48nLJbAP8KbVDxlYB/TLg+np2R24866Qp/9MN38jE14SNSMNrV+hJ
q41PHLtzloEddBsf9i+ObgicHW09laGDtOAc+s5sBf8CXwAM8m7UJarr3KtUw7IE
LlmIQ0jK5CW80Jv7wL3z4r/s8BkWh6x7FBzhMluxRMf/akHOzmxbhCKNKJQMIyv+
EHxwMZhJnbijHbDbM6HxcNT8SEO7kP6lHFQIMHqmkT11qzsXOGUIqlCKrkhUtTAE
di/ZId2JN9QPp2t6XJAngLZnYOc/V2/pv55RynDri+sQWYSUgY0uh9P6M7ZQl7cN
qJDXvTp70Fv8AsyrBO895Bjttqf3i9GqBoZDPHg6V5zkECeArT9ig+pwOM9XFpmR
5HoADXkJth5uF8VfhCrEg0FRheH+mrX1zeEJ5nA5vHfDeoXzdnfwcRRSVm8w37bV
FaIzo1pUCsViGoFBsn3evZVQt+zRGUahYLzK+UDC87VsZQH8DRJw4KzKfm6a4jjT
Wy7TCIWZET9NalDB7w8tVFTBEzWuUT23BmyPgBagFZEqCduH6p0Y7O9C4n4Lsu3x
cWHcJmTUfK0VuKVgk9KLTQLiT7jcqJ4H8xwMzCrO6hI/Gn9NERBWyoZ9xlwCArjT
+CsOsRLKiqKI1hCuN/YQUo8A3I+GvXYKRSBEzQQrJAwX1TkP+pEDf7h6K5rwZ2h8
joQO5pKycVjdaBpk6QT1+asj/g1dpH0HszksjIajBExEFm1B267VBAazp3bnAk9H
Pjf+bFNoqgSsj0B8WMuP4xl8BMHEPghLWHBdI185OVduBHxhnUr5QiGhT39XWloo
MdtabEVUdJgJgQEWve9xwzuFp5GbxSUTkVaP7IJK9I3z2pd38SQwlHWe+1qyVBsL
+ZUH2gsnYSzL5Nrlylo4Ne5MJLNE9iZVAjIwBgFvx/CEKut9bBXllmXYo2Rbf0gd
qIrHcmwcUCk6r2EEvz05Vm3UDEPiMwvxEiTcVMIuwt+CCuaT2EdF2e9jlwZPcqa9
QalKFZims99J1ZJz8jyj9JQtPGzSudC9Z2RrIT5ZGj46KaJ8AivLIoUw0LbV4SN/
xdKGj0GreCyr41wtWff/fQT7y/b4yrUYe5SxLtHVI5j5dbywbU5cvghupw8pOukb
8Vws7y2aflfCbxATtREvDjsur5uokFC0z++EpSTwa0y3d6fTOGBvnERF47m+Auet
pPowh8uGJFA+6h8D7fARYVaZhKtpK+qi5zfbxPwTWtIVY3yNPX3+0wDM8/ftLgcp
vtpg+CfwhRTgbF8flaXxxrA4KD97684WL9uB88+7UdhJ+idLNkznJ7IJh16zGBaG
wrAaXoWI7VDKib+EoTGZYDQCcEBtRyR9ad1UpRy6WQEERDFx4122ij6meRo2lo0C
h+N/ym1XFE8tCy0f9Uzs1WXJITrGSL6Reqm9FP7phNsj2msdpCfkka6BIbPj2WsO
jnBFNFE+aMmiGafFA4zWbJful9kkA4dA+c+zGAFZQ1uX+x45PIyJUtItKYlJ4jMc
hiqzFTyRi3c2/UIb7RZvL0QUMLe6e1g8mdKg0YbLK57lEBqVUtn4Xzi5DZl7zBoK
IwgnmZf+g++GozQBphp7hsqMXE0tMnpezj5HddLTmNpak6mRqyr+ZhDjNm2Ddh85
fkKQ1WGxNNEuxxUob+M+Kn0vHSZKt2T2i+dSZo40kfL75vvU0ORqM8j9H+6pVnkS
zhzrJyc0X3nrVJV6aADKblnS21z6oLIknAMpcvXD6YhZPEzS3gsgUQgWraQ63Yqs
wexvrtqObVy5F8HG6DSaN/R9pGa4ODOp5A8HdrguxO0w7dWbPjw0j+qk4qIFJfSH
7myEFRMYO/5ehCdZQo4dlyvJ7egdweDKzsfbgpdgyVr5vO2Hy80FA58fP3ZGCX9p
yOqO3RLoJ7hpaQffGVW/PSTPEvvRBzwkvCfgUUdAwCuPKShlaExiCfGrlNS80Zwc
bnY9tAKEknRui2SV72XZp/vtmURao8L21AyR2jTV3E3f8YLKDGOm+XzMHQGo2aaw
BMzys1uyPV6sJvhtuMLo+A3FHnsHtzgOJzifeW6QHeoH8lxK2I2bQiEukzSVDykp
ZQB9OEEocddtOm8klor4pkHgrQdz3m2x72VmCMBq00lquvqz6xocb8cWMt5l/xRE
GCi/Nx1KQEm3owEOFo9Cm8F4nwCvQya4mETX+mX56kGsCux+Pa+nZMTSAC44EFdD
WzxTQsakU2Gw2li8OHp80z2GJ03Xriez9e2WkXKkBhPzCwqlZY7fCwg89hq2MNEo
Lv9yAwkmBJjCQeeF2sLsksFOw7N8e1abkWr66D09814bB+pyt5YPidMcgVABtlOQ
wKGIvwwuUjiD2spJEfEA/MMc7q9eLi+ay2vAAs39PKLvmI763pgk/n056FBYvTiS
AVepYreWLjarwaLQePtSCgKFMOnKyefxz2+O6WkunsZHrjWzCV1FkfcK3FFQrq7Z
9fosYr6FZXCFhzP6Jjqlb7TkGBy6n3dRPKk3OMlEBf32Bh4B3AG0r3Qq5xknRLBJ
vcT4EXMCx+a7buL7PP8UOTBWPAsFub9V/zHVKAybIoSk1lhD2W0WlyB46v16oiTu
4Xz0jhnd7iJ8i0v1m1xFKACczlhn0dai5DW0L2t2ZyiS5Osmk6YCIi053d/bPFFB
JgP/Aj+qKTwBGX/7f4w3bN8A24vrKYyY2Km1590aaJgC+lrfHVYougs7a4JunZTN
T+2lYtdmdEn1B1I5kZPvwpH/zeqkbWlft/c4/hnrpwZogqIGRv9ZB9IoZ8aI+mHI
sgGSDgjj40TpwFg9e9sQ9cQPluDu/HLRh/DRsGLgvy8iPWWatm5W9ju26J5XTnmh
KADlcW2+daNfBofWJNjw8dRvsMTeKMZAm5muQfN0OpSbd0nGrFhQOZt/vd5er+Hd
cSn1pslggUX+7m+ZFeiYLII6j/ErVGNqAFV8AJxGP2cEYXATK9Pgt1b9UIVEWRA0
LI1sL1/XOV2Krr8aWL36JBE+/niGpNFNd9Ao9mRnQZfgqLvGATJ419wIFA379TQe
s/pyjJwXlmgTw3vqEIsh8rDYdNehJ7hkkdpMTY4mXuSPovnpNo+CluKzuSYuzM0E
B4xwhd+yLrh57w1qPp6GPFtEUf6yihV8sURtNEAVgwUFmb0BZl6TsBvHOup352br
I06vkBSwCB+5YWqKucBqOSRNm8LTFicobEFJZzIY5EFe/zmGtr4QoOguL6ghszIO
bXB7nYWM4s+GUNXGIUjnYfmj95OmSFrFL7FNjvY1hb54hRh0zqJ9upV16/IoQ5R0
cluz00W90pZ1wCfqljCZuF5uMA207Q5qkcxP9butdSrCHqMzhifOmaxeZGIbPU6L
mFofl3UgTnrRz4OVhA7e++8cYI7S1/BF2ai9KvhjuqlFmIP18pKwyhjSm3zfrrvp
GUx65UCsGmRK1z6wk+ie5bugJDTrXEqO8rSxbe6Ly45ItbMrYCw5xgnaT6qLL+AW
s1TnKYS1a3K39pTCnTk84s99hY4ZvegeZ3mQWvO6c42tvCvBNbwu/Ihbo+bCYTDZ
/zfsYzz19v68FmkoW99QQ+TrLlUweQckGHmxLCCHZBF/01B57TwBbnw9ydZHrnQX
zSXEbyih00aSqitwpSYfOAhOW0KV9+CHVFTha2mdGjAXNFd/zC3X3D+IhjtBV4Mh
rV/qxtuViTPntfiPfJl7sU/SOeylGQzRbtD/brLAS0EBYvwA9G85bW1U2NUa9jW/
Gxay5y9iq4j6g0VRh9RDTQ4qNLx5scPaSdSn9cyargxlrki0DUs1fU9JZCQZX2Tw
4lgPO/1+BXIs9wgbkInzpbLkYj0gSov/YJfg0gqhloKAzKq/nqDxZTNgSPIqktmz
kO9PO47WGumLCU5KpEZskrvz7pTiqGZsIm4KAFLG8CL3eX4Zx8N9LSBG70m+AGJY
Ah3QsNOfMc6U7RBWoQjodR5J2vaYNimn6FMYOAWykiH/iPEvI5esQG/60buqZG9o
oRqO682shTcl7khX0akUJx11YPkxkNGJOJLXLyH4pfp3uLxOA2XdlxmfloMW703G
eT9Whbete5n1aJkJnfJwaYX/7QojyCr4f/V2Z4eGdfCZmbkXwUoBiwSbjG8K/gWJ
CoU6Qe3Y4Zi9G6Wnk/TjdQra0TVo3ud1hi020t6pWZGvvLqsCqdL9e8me48LVyLM
LZ6Bl+xWotY6loeXFLA3bH1wFFBiaurd/8zXE3cyKieKOAT6Q0RQGC17fql9dlPV
yFkKtv/PiDiQmSxu2TJB1e2L1wQo2pmjFFaPVEQZRBHDPZD6Qnb+qgtmsfSPeClY
Ix5bCuD6PwnfLo9PsvN1c3PSMWEnyW0bgNPkEqa+BU60LMZiX681lPvTmAgKZ/Vk
2WzaCxqj+5+LMnr7vU7fDKEvmzasHYwruX+96zYQN9aWh/K4+OfAxqCzx0oNvjOc
e+deSAJuTh5f62W7HeaHoqFGh71ATOJeB2Je3X1cFo4jgADqfn09HwwecImbttNc
3qY1i50DVuGTRSuf5uW6Mry+fX3WKcKJ2eKeMGxFH6XqonpqAz18hz6W3POU79j5
fo6A9Bnmm9aA5v53HuSnOJriSsITqPTEEfBGfbxpuoirGr0ECmFFWDJrHwQxS08l
CswjIAYqhhQrj1s37bQFxgXknwueH9jyUgF2oJyshSfa0Tpl5z5siu/mxa9AjyKN
9e0ovy0k23urGJjRT3ZVZ+ce8TTCOXkRReNLXa6/szO4NmqcovCqUb+3ZYYAFgWQ
dIflN1PAvJgcYHDKyAAWy0qgpo2DEtucTr0As4cun+BPwXbgKyOcDWCoDZgocSew
5IrzfzCDGTHkwWhV3043PpslSMTJu+gE8DJ6j7FQ/mQYaWu1emBQpwJJp47R304s
NWf0bc4QhaGgnanXzJKTnEh4Npt+0TSbfWajEgIuV01SX+22+dDejqXDH81znruR
i1Y7A1bh1d/pB7Z+B75c6q/UchsF6m8Tam51wBU8UKbloFXBpRdOO/nrRKh6Es31
DsseYPwgVZ365haK04449SlWQqjInba5j29Gz9OxuvVn1ySJmbAIi6cIAkmfskA/
BQKlFDKpQNDq4sb8YKUBakIS90xOcSfBGRQuMzQWa2I01jr1fWdHnRZsBZ0vK/hN
xr9gkl71pVNdb5LECwlAH1yO9rfikxSCMR5yNLwJobvzIcRTIJUQ/rd+08Iu4y7o
Zql6sRhyGlp4jc4/DWu9OKvzyk6SBIZ/TrvNgdZyzpedpNIS5/tJ366UuBxzP0IB
YhvgMgsaifNDWdxDjSqEhmaJZH/tCRpRTmpXchj4Zqr7Lw3paqr3Sw35d0UHvFgx
IWma+VstpFvWuxQvOSMGT19o4VZC6+AszrWU6NJhrfA6xzJ/dlbEh51HdkIpap4J
Fs8ygRLu+4T/9jRrhg5V7enybTCqlg2uh7yHxQ/W0kNaraoGG2fLHEQUEaE91Fdy
Kb3p5m/vmLmxXagk9sDu4s0W/N3fC3IltmhI2IbUERyK1LKIFRH9KdLFVX9njI10
JO8ixj8AwjjInyLdE4NTKzw/ccl/llQsRlGZMFZNBRDn54RuzUVIacfdjYSnKvRW
tbl6u+ISst1Fg13epnoZjYpalPLeIU1eZwk3xTFDF/91egn88XZtJX3Jrx1SFpEn
vaSE+mtERczcYufvUnkqeLXlDvCpxENy3nmUWvPvvUMOMAMqn4Qiz8xWKsL0tiQ4
EcF1fCj5epqSSnTbMRJp9Dh9y5Z6Ie0tE8Cv5hS4MUimu+QhjPJgu+KCLSf4G64D
FZyYmZgQwSjFo0pHkN77VEle8DF3MoIGsCVsAY2v0lLUbGgEzYi9TcnPVnMy4bmZ
labJw0nWvfYZgOSmG1McAkewivV6VKjc5xdEvco4fO5p0TWN7d7Jx0NbLtEGmWru
lJtcFwDMdXuo9OyC9y+KpTXA2X/NpANnrk3tUPWuUmQP/LMz3csR4tJH7t8+bbHW
VlzjbnAm8zVLJpA4yP+33bQS89XOUtO/5GOkjAiiONx6KCwlD3NC6S/pRx/Zyzys
aMV5wDhhFuJqSt5theatYvHxpiW4QDoo7j0z4XYnPnc1u0c0G9XJ+QsJWw+tYdMC
vKfzHU0zphBKzkWC7OtLL6TAR/QAeZOZ5FGnyGvEWtqbC9SXWnwYVOJqPEnwpmnm
Bw0nAC9w2SsNK1nGLFSOPcvoVtCiqkjW2lRqCuv/wt7KfOaKBicwr1D45cjP6rXB
NUxAJhDbcQHZZdQ3Xptg05spsemLftI1gBuwUafkHyS4Q2nI2WY18lTS93LtbNLY
LuGnucTtPQhj7GJWRFjI9EuKfncIJvrTJgeA3rLjH/TCQr3uA+ka63a8qXvcXO/5
agpkj3DaTZmxnT+5P72gmShJ4yaj6EHycJYEsM+GDruFw5Qz89aG9L7muIiCtUW+
/WNmP1a+68dCTFZzppauMS4OvLJmyuND3ps/qa0M21mWGECC2nyAlnMs+x7k974w
nHUg7SkeH0A/hbob8WMBKx2txxmyXuNHiCydP69aHDD3oUTfG0i5N1IiAsfhjQNc
tDsVCzsOVtz09bepusxzSSLrDzyBkBtDf8dkl1WFLFMjOifgZtFPymAwR+DxymOl
8maL3ey5+FSUfoFWsAn+Khx+VXJkHexLjbbTAyiBecrrhmb97I2WyXkS6NaNOr+B
c8v+/YlyXg7lRs+pLgxJSExlFTZ+iy16zhN0PBAxqJqrmUV8Ciy57SCROry2Kpsb
6seLGymibjlBwlx7/ht5zOvdddZjTU3C/gVS4ECrZ/+Npf0ooXx9XtDxASgN6rGt
19FBQYFji7Xd+EIc7qQhVoxjzVkDULmZ05MxUpwx5j3uObpoKU4e4AjXCHPzdNJD
cYepNRfur68IKeY0OrXkIR0yU8INlJgNa/A917BNdJaCV1AkGqvUXnmZZQUaUuKO
Zp5SiDU1/UwX9Vq5pq6VDJsNnKelS3adYhtnSqjMFsTef6xSx+CZjfwi6PidgUqY
DUbqdiuSWxne2tVZmek8taZqxL4Joqcw1KjsbVDZGeLXsIZIf48IaGfSm9bli9eE
D9PMK343Zpriph/zCCXKBw5rEIdNuNb6KMW2+r1PI+uzeJIzanFOMzvXW7mTBSth
7DfEjRupGTn6u/CZzBxwgaaDYCcRhmLx9fUEKSS4IGtbzMbMYSiP6M72G6rCFLUz
DV8rYEHZFy4ikxkigPZ+uxQK0OJDCVQxN0FtOM8O6SYc8IXIR71JXoDuh9Ad3vyx
aeqDAGljQBzs6AKY1axGExAlHJnx3ah3Nbyv7zWp7ub1m4ehKk3J6RSl1w+xOg4L
aljJs5bYzE6f82oCefb1VFXHm8MrsyK8k2AqVWeac460FwzAFfKxJ2iditatjZOT
ANF4M9ltJJE4ZAEJrElcZVYgO6kjJ7pOzbb4zr5nNHkR+W8Fg04ONdTH3w02OKM6
xoy8NvtbrKSJhmvBUiis1FokAwg6aI2hnTtJLGy1me/2Ys0AwDgkrzYDpxdsEINQ
xo2sLzv04ryxEU0hg2sIoHnZvwI9cPN3luGgKEM0g/unp9CFDc1FWW+Zd02l3gO9
v4v3Gm1jlYDmBJTZtB40tjJ3WkUvjFjYH30l3GRzVNYVBI1I4H8dA9GwhF9c/VUf
rNz7m1hQIiYjKrOLywNC1+Aqj9G99e5Lr2vLojNOruZo1UG8uWCI862mETQE4kvw
VbGIkl/u6NrR3x5eghmUC1gJoeIShlcnTDSj11xvQnDh+VcYqREwiUQUE2LMMSrY
TQfnzvLS5FUrU0sAnb5zUgTXSEc/WqEd/BQToVYE2uKik6cwZ+d7XmibDtebMO/H
CXk/ne4JxukcsJYRMHMbhVJjVKHU3YoAzPnGkUwCEs8vzHmXpVAM4K7OoxichVNs
ms7QGWucLjNShGobLzU8o1zUTvdOiH1zx09Z3ylNrQninl/OzhCJjILiIC+KAzNA
8WOAqc/YnYilyI+4rKMd+7uhiOHjwciJwLhY7zfnG5+6yFpsqvAipMIypiKUwUjV
MpH+rDjoukpFthD8tA2L7leoz5snKfrAcscQYetdCyxmnyb5VP5dYjDSSGutpR0A
dW9jHMNadhYTa1jyblOJW96t9lee6buz4VaKNEMEeQXCc2fo/w08VhSNBtc/XMkn
yfd6Qqd31//JqsbaqwVIbps7AH/Ip1Y5XWjtY9Qfx88S+Hut+KreRa66kLk+CYwW
HlBYG8DtPYXdd4TGb+2NA4dOfDkZNEACjTOXj13duvl/QZaEAV3LOvnBNlWJb2eO
2SUwiyhJZy5e7Exy3x8lY0/HA9QkAoxGRD4g+GQXxN2kEB+nsGi8h+IvVTFRLt7+
kUYlWX7ubkPXZ4x9OEKwK7avMbNqy5AEomQDP2HLosfWYt6pXANDau1R6DXM06N5
P8mVNiwDKmwNFvg/v0PIyZR6IzRKap4GOjKQnCHtUESwV0+ho/+IxBVOu8VS0CH8
0WqvIUryNhliSjx2zgd6a9mKzGOReVTD1iDuajc2uVHWzlmWvp5hL6+adjvLo/3n
Z9Df7xbnNngAEW8Z0jtT2+0baiXmJg5QUB4mxrFIuM/SwEift0TE0yMRMZqaAReL
vN4pcriwrFmsN9kHgPoNF9uRy6WxoBREiKYdSgUbVE9vZUN/Xe5pNyO2SKjqE8kg
PEmc8rqZag+HCJzVMAGT/LgnA0jn7y8kFS5h7ZiKnTdfNi4tYWOeaOVHb8D5qF+p
rE1nEzUXCMQikykURmbFpda6FpwB7jvnVzxTX06+o1Za7Rd4I/Ht0QxpukwrXaqq
Z8VUiK+TbqjCmwsy0umxmYv8THcuKgXUaF2a+v81cpgx0uNjZ2FPxgbaGKC4LLio
t6UsRcOuPrFy1UYDqU9oxT0TiyWttRZhm3bUyYFhf5HfkasuptddL0iaaYwzf61a
YJX7LIFYT8AhZLXhu1pisw0wm+5o0Q3Bqo94Ek2PnnQ1v7SAQVCDYOi7kzkNU7kz
8+hAcL610U8gLoi5zPajzxf54nLB0K6sSXdC+b2x3mihyeZOu5URy4qzTj+HxhLu
reh8mgYzDyqe5uxePDqn0e6rvmmlLkTn5LlMaT5bcQqnlz7C20zbbm7MeCFfu2oy
sOoiINiPqzGHyNox7/Kr4HDqDP4vR3JazZdH2608uzduLbWalnmGVcbX7gNwealf
c2OvrpMG/NmXf++onZa1ML1J6mJ4m1GaXstuCUYTyVqYqgbQMaDxomZrY85zWP9U
9nAnyUe6jzNw6G0g4Y1Zn7ISmxwAtBJgkdVBejkgGWQqCvZ18L1GnOQHijwUH0Hh
LTOD3K9Z/k4BXOoR1OdF3oh4wQXJKUi7Mz9ytqL3YMKaNVxvUHaLLGTzUu0/81lD
30wa15Q8mlOKDX11d8J4+gccYJqzqm4Df6dbDT7Zdr+OOuYh0xb89UGY8FBoIISJ
qg09WxOcQcb4QnaJ1/5JQiV3uAsPp002Hw3prPOU9RDe12ZBA+LAqcT8tDlKCa/S
jzO2XX6W5suOaLtlSAJfyEUM3gMCuvlbgrMQ95roZSz1F/oskvepzIZqlrh2vg5H
fnlvWm+7/btFIljM9Ng52cAcLE8+Mlvef/HvOrr4sGPsFHgrZ7NavG9njrDY1Ri/
nx9WZ5uNyDjS3D37pWtL7VS9QtFy3awKiPZ2k9kgg/Q5ntryimrKIw0dzFHjdtJD
Kf0TyjYloLanAC6XVkDNpnMLr36ocMVbH0QZYR0O4M7Xj5NLYHXm5MVIjR/UtRVj
ZFg5bO13tGs/TtX+/+iwLUbXFFwT53qUp8u+8p3wm/qQrrkENJMatn4Pqyi5QA6o
CwSNS4t5nuDbJ9SdaSIKMvERp3JIn0HrwPHDp/P5Lzc0RBIu/aX/uED5jXCAat/p
sxLK4aOxDENPJn5tA6Tn/hbWdsPhQFUboe6oGRjEsDwZB/PH7pzkIk0r0rhgJD/q
XTwfsljrc3ALs3GSBBaxaPtfA9wIBwt7WieHf09qdBWCXVC2dFtEZlwn6QX2tLY0
UIRjCrwiFTgTtgRHIL4X49vEY902iBb/th/MiLB/tOknzu31p+shw1FmhgSp3Qy7
IP6KosJlc15EHY0YlBi5Xtvg3/yDz8cZ2Pz7xZ4deuVvK7o9xl4XWwT6lPaPc4i7
rUdWLhE9JwLTf/i/il3YOF4DdMUSQgJiRPfNMwKrVjfv7LWy1Vz8dQf3OU/Z7t5F
bK+ixNliYr76tfQMEGHSkrpH9StGy3LbRd2ss48CXErvuRpgWniThR1dR9k9y4gI
jepIMYCK980WWLHINxcpGezwmApMBlCEbYxJQigsfgy4ngoL4yNVOHY2gjB+aoFS
ADUpVc+ANqEE4sH4wlOhAxhpC1plbwGLRJyn8RIWmWXvuSspoBb2fiodE6HHu7dU
IZQJwRIBTNlzy8/WOqQYp8Na6i+87HHgTbg9g6UaKOG5yR79Z2hsff7AsDxyrr5a
Y4TzKLD418JgjSp57gFHYO/GDXepCdAZqODRXyQAw4ya/aHiXs+QqI9LSPv6oZyJ
zytYWI5PsYJBUsgubYJO6hz8IFmaV9+Bh2VNX+8Fy5BgJbWtZMFJzhZAlkT1wQTJ
bBIT+RGNfqby5GjLKr/v3dKbf4ntevMthV97ZDIOvBHdAcemisu7W6DHHvBtaC6Q
7XrAGNGmZcdJFhtC022g2HmJd9qF8b5ULMX9ffCMsFENfiXxYD2pdM964Qjvp5Hs
hKccSWan1CAntAsPki1hPlKOad01CFMzLlXvt1pnNVQTVg0ufzmeXaE6nZWxS47B
d2rv8i4ptzcTZs+diWkr0jronZ0l9AYaAVpBolBRTKm7DY9CaGIjhlbTxk8hC/WT
TQUZlOfQRCEgPzEmMFOu+H8GC337rDtLCPJ07q1UxqNXcxPISktfBErl+7a+I6j5
IMAfdvBU8A9Vp+HgqaDnW8NDQhzBNzeiZJ+gzVPMdFCC2QxsfKmcujXkCr7sJLMq
dQLnUjmMuyiQbXTcNXQM/7xpaHjEgZBKWcqbD4Pvi0OmPrZDXmOUOVgUx/pS41Ar
mybLuXwfd9JlGJR7v+r72z2frucBB5wJnABK1+FkDqYhvpmQQJf85Ln1HGdR8Tbu
MPn9waMH6DBFwh1wvMUyilGXK+HTjBAeuMWzD8+v7ZWwx/C04qPmT2EHMcteprJP
UPfncTKYnBspTmJ4HbghdYf8yGyy3kuHBpvBMQ03HUZQEGrE51vV8xZL4i5QEXto
kKnAAZ8Q3LmFAjXlfn9yaAtqEbtROpDwrYGMiXcQ7ButOxcKlV8DdrUg1dkrb1oP
jcX5mxMC5a6sNZ4lre+xO8tytwZXPxO9FDhrPjI/W6Am/aY+7GA2/iV4EF3DBDMa
b8ARi/lK6aUMdjtSUxfVHkZGpkjrFdvLPNLxRGcQReTC62bFHjAXClq1FU4XJ1d7
Nnb7gzTk9H+mh966boxbKbQ3a19S77pXa3jyqqjZPyNCrVb8B9dS12PGmKSXMtgW

//pragma protect end_data_block
//pragma protect digest_block
2eB8uQIv57AwaiSq/+hgbr8BCIM=
//pragma protect end_digest_block
//pragma protect end_protected
