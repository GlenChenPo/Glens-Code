//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
EiaJDhBRuaZYOYxziZDV1Ymp8HLNnWcK0vMDBlXkilKOQrORkBthzb7wC3AE/JAi
kSYqO5KICW+hExDN7Lz2QFaxH6Cnar9QhKu6u96iKuWJ2NjWHEUSbgUdxPOP780+
MteW0zUJr58uNXTmX8LeU4LQaHCf9O8MlTlgUpWfv7eL2gU7aup7Vw==
//pragma protect end_key_block
//pragma protect digest_block
dGsG7weH5VC2ZUcN0MmeuQg0i1g=
//pragma protect end_digest_block
//pragma protect data_block
n8PO3O7dE+YZMID7vizGZ8GE8wq+G5KUUvJsx2Fb3RjRf0yWfN8/ioxxPJIAtOsL
AnNILgtt+LVGCXEBFFExNAmZ2qxnyHQ2WAjuH5nCi7sI8emK/nFHfN9AYsKtifWs
eQ0ox8vReiEOAsdVk+h2JwwboG1yv7G2TVlO0u8ZEXAlT/JyvT58hzIfgA/Bfsr2
k93b8xDLkHROVxsjsiETjS27Nf4cY3/rdqo0AuX077WFuD0djH4N7rrzAJE6BF4r
R0b/5EkI6ueTlzkyfFzvBND5QKElfN7rHfcrN23FtnIg2gzsVl6Ap1iV6w90n5Rx
DS0a8d9snDf6zS8LWmL4WQ==
//pragma protect end_data_block
//pragma protect digest_block
rNxY4y9bJq7CWl3GwTA7ihI1Ks8=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IZ7janS0OghugJ6JFn8tlnMPtNjBevQ1ekQCjrW/s8f3R0X35aBxcDbMS1hZBxbb
kGaj8Xg//JUQ2NCKL/r9KTt6yi2OAb0OXC1qvj8iW9eanTMFfmOQC6T7vq/2srpa
Tdf6+QN0es5X6CbiXzmWPEf4+XLs00aqNmmyG1Yyv5z8K0QiTLcX8g==
//pragma protect end_key_block
//pragma protect digest_block
75iDT90qP88mt+f3ox9f/4U1kFI=
//pragma protect end_digest_block
//pragma protect data_block
p9FgdxOMEqC+SITqPLXezC3a6zc3M2ELHsq5FRHoDp/8e/UJOtB1j/01puhnwdfX
g4gzKsvb2HmbadJum7zO2RrsugJRS/j7KrgLFklWRmMfTufHzs4iYa3foxYrTyO/
zpmYmArS6QEaHzLthGFShsgrPjqqqMa9Ju0qC5XRNfz8qIqjJH3Qrgm/aWEnGzZB
udDZDSbflk4vZx2ixitjKY3IN71nzwwm9mog9X48HE+eVUK3N9G66YxklZbIF0Zp
4HOJuw+EyxY+EEuh3jfezzGUzPhDz6oq3rjh1tKvl66NJWXPBjvNDT2CM6mXhs0I
b0Dl8TA9rFCTqLSjCnBUlw==
//pragma protect end_data_block
//pragma protect digest_block
JsKImzevSCWrrK9YCnFpDhCIy7A=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DYKHHLROCK4577vO470vMqDGD0TAmcRzMYmMlOaP/e0Rv19RcKKck5HnjDUKLUXM
P1yd8rTd2uCaFfB8xbWZBJq7kn/WQ5Z21fly001Z3DTtnsmx9kVGeqqrlKGKFqV5
IPifNLShb/qJa0q4Q+JGd2mF9d94ZQblgqIpRswDDxmba4JdY6mmZQ==
//pragma protect end_key_block
//pragma protect digest_block
ahaZLtPpjTLAB3kAaNaTvkDyqSY=
//pragma protect end_digest_block
//pragma protect data_block
LgJX1wFHmILONddnCYJV0UP7iQ2tYLEKq/PVSXXH4pIGW5tO3p2eEjyyUvxnQGbp
U+LB/pJqNzOIR6BTTgRYMs+2341tT7RCVWGpmS3+YZf8LHZ4jSZccRMaElsvhEYP
3gM739onAc/5NGo9fHEXDChzivvyONaPwR4hrrKUhp4rI1ptCocxE4mG/GCCuqgs
TrcaN3JMoVu2xTwaTdISkFCg1EHkwpPGoxF24p2G12G1gqLFHyoQtc1C4NdSyyat
9UtKBEkgt4GdUHR5vLjQ2o08zBa2WeItoI67E1al61aw8RW6jMI/TAGzXV0PffrF
cQMSmoBiBasJZT2qf+a+3PXtaEFSvPOYBIz0UKnD6S+tvxhyLl1yrmTiq09OmFWm
P6tyD4xkcWqCwU3lZsJ6aIrC6qASvMQGfw/T8LpcX36T4TiVTcJeKJSdnowaiNdD
YKZ38ptUXLN82eHbgsXuPtfmsQO+0WMhrrDtahli60+24MNn5CV9ybejsw8oVdyr
87Mh+Jk+jz4xnw4q1aZtGsYOGvloVbG3lwzZOp9jzTrql2dSSQBz5hfY6tLt3Rsy
DEr0wgQ+RoChOa65/ZsijOXCJYZdPHZt1Up0EhNd2Y06YbANzpd4IO+NLAPig2Sw
mGzzkUAvJXgMgHXFB3crOw6d9upDf2FGwLldX6TkUl+uyAalMiLa6M+NKjEOQbQN
El1a6L2bz0k+JGkYmM05yPG2rIpbVergDowG15D7TFt9IxWN87XcaLCQhlFpLx9P
54ilSXDZSV3IsTOQWK2O3T1j/aT8qtYlWKnYF3lsopAdebuyGjn+/3vrA99MU/Cq
gdq9rcTyaEYWlOpfeVn+fHN9x0kU2b2GAcFyXCAx5WKXy9FV8sV+wvcNXV4emobd
urouqwpb9mgQy/dGsbFQGWqwlps5Wc7z6z00TLILnH7X9dRvvfRinOLGxoIgii9y
ZldHThQmK+IjF9OVWp3x6dc8p3YZQ1iJ7rc8IZyFiA5EMdmDLu7L5q+coAE4TDag
gtDFPYjHmjifvaBVnyHZWyP/1JslH1EmCiCrfVo8F2YlefY1MVg1aY/TJBdBwdcr
ri9wZDJAO45t/UDLorI34AWuX5KymrB3EcASoQSg75x3k7iGyb1+ZSpSMkq1nFqP
DV5lXDUdg+KATSKNyfWWR4c5FCttbAb8naB8wH553WMbzjXNfUFtdYXmzJs+h2pf
wlvpIwYt1xApoldNO+zuiLPF90knWXv+mKRhjSk0YxF/KQOc5nT+yq5lwfhrrspr
C2Rto2Q60I3tgH9gBPfmXI0+ZmmpCd/1tk9W3y1uR7hq3zSnjdXlIMJhjlb7tIK7
ogmNj2mAQT3VSBJs16O3viRjudNP8FebSvFeusRkLJzFOe9G6f+Y0lX4ZdnNeexf
Of/NM3ESetjN0n69m2GPEredG46yxbIKs0NvuVFk1ameyIeyhrGg0md3UivE8BIS
9bCAHHj3les2lkW/jqmQvPW8W/VJKfBSKiXuEnIiw0lt+XEJxQSJkUAR/rUKO3N9
F72uGbq13x83I9beVZrKWS4LP9U1NkVTq+/AFBm5ijt0ffG0LQ5dACfvM+VSKxsU
PQISiJmmUTczTjNXWdDI/BU9HXre56OyiMv4MzsI9MkGfVI2wNv6makvBGk+c4GF
bS2PhEVeQa8CSEUgdquZX6DVmafyeE62wDqD3xuTVK5eMvBLp+jkc4Wxpt+F44P3
R47cfhbR4VsZmhWpDd40BESLc6e560fzlQcgvmF2zeUlNqzf1jvNRAGKKCjTCQrk
wWr1NoL2el/9CxZ3EV7qhI/9dINEltsjLMhzsFhh58iU700LbXmlWhuEpEz1oQ2j
CFSuRjKHyZKBLjxQXmu4WRdGi30zYCURHQwybUPVYiXpRcN7QjvIScu4jPVTpjf8
+Hm+EFZKsrFh5jdYtKSMt9R98EJE7f+dcr2dweLGAc2wsusWQyO9BhY+p6NDbODh
sQSiE/Aub0I/OA1o8f0G7hEc6fACC5trGqsDo8LgxiWTqt1R74GzMU/95MpCJy4W
GW4N5qUEAlgVCl30dsUU0dR08x4jKwx2dUr5Knyl7/eJ//YXKZBONeqwSh4f7+4a
LeLVxqKfzIXCUutBuLvp11ZCBDOq87Q1P5odbzS+GdcaaCRAXZFf0SEUuYgN6qy/
oPpVNrFkubOW8qx+tKCKGOZ3Lb6Sivu/5PYnPcjZdpBRFAxFYvdBB63YcCNAW5Y4
aLmI1esf4aSJKUtCV3KzzB+Hd2km70pTL25AW0QkdbiiT7eohUyPoPxFNGH8tRio
BHXENSzSwekwOaPjuagLpLBIoB5wW3L6SgFeomhXI/x0KGv+xVYV12e4whd+yPCM
xbm515tbRxcXsh6koQLQtF6EXvI+aV53oPQQRDqDXjgoiaKxuzqvqeFfU/TE8yXW
yKC2GAAfl5TcFOkVAKq8p3m98WdG1Fo2IwlDbYQjnozcNKEwhH0OGc3zEovVAZoe
tt9lgpnWR65SXvEpLdUT89X2lcAGwI0ny4GulAeyR1Fh+mtVmOuNVU+XSch80ox2
Ip2Vsg2i6lsCTpI6gH8/6ogSL/dDDyYbUpEPTYXXS4av+1CIIFFob4ZJHOI+dYjn
D1MrxHF+VFaF0CUY3acsD3QwcfR5rx0h85zLmWPa9ucNzPZXDch2QEYB/AgjXTKT
ARgPuPfjbxD9GrQerjL1w1R/rGAwhAbf/cbcLQ81PWOZTLCk/xeFAK7iIbXDBHOi
Mz9tCYVVFny703Hgrs0Uv6Bm5fdtlSKS91aG1tsSmk3fE1mefDCKVSUxgqtegNhJ
7PpT51cEchMadRBpPlFXD8Crfn2mwekCVgXNryKb56YJ0qYJ7s1xtU0dIMJKcB1t
smcVRjnwd8gFmWSCzR+ju3iIUqd3tR8FjthOMVpGzUv2vZFDmxtZtahZFfo0+3L1
3hEX4qEB930EnT8riV2MBIqrFOyGoOdKskGIEMLxYXiKbetEUiS24gjY0V+aN7zf
yd6Gx8p5K7h+Yomxso5AsEqb7Rhp0wkbkecEQNBFIQBfeYyTnjSblpv14Rj8lwpS
hvSQxhTeTCDbq/ixtWQlzc4Mr/T6SOP07+VC+1mvSSPwwlDLtcT00CwrzwFwOWUs
/ekEeTtljvckfEjuHVFAmhvZoBDDYStrDBAg/dPK2/FgBOsmLAsgxsou1NsjSRol
J/2KA7dfuu0HJDvQdcHkBJ3WrTp0xemJW+nTzkqFlBTyGW3jOzuoRVAX3gFLJVFc
IHDFZFURV6Afhdl7/IowcbaR26RKiuGS+AE9GpgO2fC2fLHe8yjkqq45NDVhT9yv
WGVXtwfQFwlXuHQ5c75wPgJAUC8zgyC5wFomt/3sk1tTsx57kp2i4ziSwYx4tcsh
YqWWc0IC+D1/GreRvInmlgBdN24TE4iI1/rRJBmr1mKPYSMdngdfWLFw6zuOaMhR
QCAjj5Psn6Vx0wrPQ6CVP3aocATaUnSMKDVK1YnWfItKphFgzmLKLXAOy9FjIQDN
tircFAxIk0Huips2tYPV28NutAqx0luE1FS6s/2tQcLX//NxdCdMlsRdhM1/6Hq6
QLrl5AbIpFcD7kdIbKRWvbLVXme+mPbgZj7X+KlVGI4ugSNfRaY6tOwEquGWTUNr
HdwRb4aZLJ0l6//hA+dkc4gtDL6Ay41kuy4VE66/8OEpmmxLbYyItdf2a9C3VDnM
FQBYTFBqm90oiP1yrETm/P6OnZIKtpRe/mbcSDPNbVWsetqi/ZyaTOx0ZLuD3Cmn
iT5bwwuoMtBheZVHaDKlW5LGLYqwqf/4kKCSdHIey7ydsxN3f1PWLbxseibMu9r4
8XO08P4YjSKfXA7prnKmXxrVXZWTG8qjgXqB5ndXGO3CgNrvi3jzLthnHDYdtv0T
wyn9UGozhqZ1mop3vZiDIzmt5qd3bkJHbIFPxCxii0AQjd3pxeS1m3/XV3xu0b7p
D7PKykWvnoScs3md2vIhQbrgW3Mf27DuKuu00d5kE8xNfG30fAxTJq6gSzNl87OF
6b8E75OPtuvwmHpkIK2Q9tw2sLadIPeO7AH+rRFRTXgKwF32WVx5zj/OMy8OuYP4
d7qUNQIC4/alGG2jYqNsZ0+NhECjyXkGDsPpCakVTt2m8k5FXKjbEVzTmJg/mNX9
MdFjuJcbUI24Hiq34RO1npjTsufkS9sSJ0CwdeoovT4vPumMm7PX+NwykPxr+85+
9sWFQl69lUr7adTVSYeVaSxhB/5pMn2Do3me27o1j3qhHo9D7sY/XvaYWrK6f00p
Rbfx7Sx2p81AXYAnQJvgOeoexxsyG31sxqgA8ta/wV524iScv7oSeh7lfzqSNbrz
ZnxaKiEpINTjVwDkbTbc+k369Dy/VUwB5aiDc7urCHd8Puxem6qSJ6KUuzcvqWVH
JhBVJv1RXix140IVFEHRl8gf8kE2jwY8vIR1ppDJmx1n83AfpJjYagxoL5fcaWsI
BSAfkVFdWaF4i0f7H4oX2sH9DY2JVFibuxYLoWYJRryM8/OAwhMoEidR0OPcZ8vi
ne+KqJCAm9OyMjz/ADOHN5Ys3hPiNjoNwWs83wc8/W4WyaRHUA3aZbJP/nGkofNY
+UvoXJWOFgs5dbfmQIIitQFeQStgmZHl3FUmmtrU/lDMqVuZOBb1A7n3UooScT/n
DlPoJ7+LH5jOFXw+7ONbK6ALBJjXO5hm+8sSYIN4NBEyHjipInML+Fs1IfUomEPE
jvaVo1GlUQWPcEMC5TybwbBxWoEl4TMThSQyusEwwcNEz1fIpG7dzkjrVcTBqxGS
GNq40C7mR4K47odrcIseMmIwaKS3E8sOSVyZZz1bdVktsvOyL27me9/7WVbVB9ti
+lm5ttPkDzLNncmD/ZhZ+q8g/sQC2DB7ACcNq9WSfG0zUHykHCGxAczEttsF5R+n
HaFUh//3zXEPEhQQitmH2mSBB5YJkXDlsQIut5+YqPQX4FkJq9BI1EtAODcVPLNK
Td3wZS9svuFWkdf4bWEqR2puLum/3kMqhptltyTFEeYP6chAfWSXWKmv5LGRgviP
e4S5SOPO6J1jewnDFAezvZcI1IUR+LctQ8IljKeLTlD8RbAGpyCaagr/5jzw7kRd
VNUI1QDiK/weFhHD+PrEEFE6Q2M8rEgj6OwELl32G/hzgUeOj6EZnBpfAcUnpYYH
luxL7IOKcDamlmfQyNDq1+Jy68lGg8qI1bsLdroeBxE1D1ksG6qdoRyX0iHmmrLY
gxC8wnToMVPRbaQ/0RHuYb10gY/11CPeBAorXu+gn5T2d1gBMYoOfgmdJ6FiVj6W
v0aJdrxazL7jOiXgRdk+Nqo8cd+hBGuTS7AP6Dg6Qfj6K75iwRIzJku7LWNVLapc
73zcUDc3CIAL8bb07PzfMesZmk4/lXdjUz/xoGYXF7BYbuOaiK7n9c1Wat35ZYQV
FCci4+WfkC35zJP8BR+ZwgSVtjsT0vu7pTKKtaDhEiALv5YvY4ZAX3udo4n73W5X
T7EuQMpbP1F8HuBKA1XSodkPgHJbbIv7mmtPzap/F6lNBn9B5RCGsBnyUykdfqg9
nnvqvS/lCF8Hlg86+2s3xUKrb8/5gEiOePOIE9RfWa27ycXBvFpwXjAlgoRfom8z
7c/e/+fyXYw5dyvVGwSvNigQSDXe0rzIRleeyYZvPfiNOSfgvCoDcIczHBunCSPK
pjyoEuIvIRvkNMC8ayhv6xbFVGOcLsgn/H/smRW60VZAyBWp6wOiFYCxFgtR6+z1
Zzgl/zAbDfIvEH3ldFeU7JjPgnz45hvs07u2pk1y7NomaiDp/xG36zyi4hLU29g5
dU+w4JRfXlzccyHfZkayuR7/IPJzeXNSpqKRo9qvcpySjyRmk08WoX5igy89M8A5
uerhT/1Drfp6cRY4FJtioRF+QFi2lCRtEy6UscQD8K4hbsfw2tjzPbR5R+RjWKJW
+rPqthwEkSH9bw1nPwHJjMKXyTyooj69/9QOMRKhp5ffFp/LQJQ0K4HOgowHgUcT
w2hqEnb2fEOcoXwNOYYwZbiovJnqcerx/xsreb+Ayu5WuqJp2YZ6RrOql3GWzhMa
xokSLg9fcD4wfz2Bcrdg3OtAm/Gy/1DspoMklQ3LojaN9mhDh2k5GehEOObFN4yA
m9p216NeU5HRtObG0MNALTvWl8Z/bRdzF/Ce2pj5lcZN234/KcYoev3Lntbt6DX1
gPYs3p4iUOcgcGYxRQBfR5l/AU5r0HJYWHR/m+dRBZvZLavE/KOa8As9JBjwgXpR
cu5Bm1j63D0/5R3IyzhAwiIRjsZ7L7ATrLgouwLunkFulpdQetN9tJ1+98ByiMo1
JsfNeC5QLELpxVWvsHT/1g7O3IKy6YASeELJEVC63zPOxZuj3KVwUwpv8mv3TOYe
W/GH6kcOCLYn3MBoHQ2BNCjXUyDpugvnQ423y/SfK8Ur0tpM2mN0UaHHx5SrVkyB
VOa/8iM0Uc6dipQEuu2U64ghREMpJX7xtRkzrZ7PKL/wO9KrNJfkrjM03MW00KWJ
gH01xM7Ji9bgfOzNp1gs/GD6VgAkhXbTZcNkdrkdRWZOYg9NNkwBg3AJ8uxxbt2T
N+B06ZgQ0A+XD5U1HkfsIoeaG3rvYXbXkK3IBixAzur6Q+xShBVx6McKzyUxMIb/
hasz4DhMb/2+Lew9SlzkYitHxXVMq1n6xAWnmBd+8oveC5KqG91/a7Tu26/31Cls
kG8WMkwg4T1/0uNVBCJQH7vJ9Kd/PZxty8jWFPeeXq/J4msHkmIUaoJZtyJkE9y5
W4o+1zm94rQZl5ch49kIAt2ceaANoOH37tpj5m5UDCKmr3Jc8ipMkHaaKG5Ex0+x
08wHBwOScxYdDLEQGRyDLvqsucWX0r6I1maJ7zdCgSU1ggqso7TbY/Lecj/W6xQv
PEKR7jsooNAcdD4KRb1ed7wAP9gAvOECO8CZpFSNbDXrJze4wAK0AmcYeetcxyAA
lzxdPx0OuTpzg10eSfLg7CUSIsuHov6QMegzUGBYZVOv+AfbZP1DjYLZrFYNOTXT
/uJl2s6KzdjlRDu058W8BHvyv9OhGIyJh8hG3F9sIHjFb0x4IE8H7imtoYIU2QZt
RHH4VAazno16YLL86wKjPk5bXFBiqkZR5z53Ili08KoMhlUk/OU6fMVT54v/JMwy
qfDC9j3PId+SY2oMCnjvP+1THieAgJyEcXu3kVzT3bIyvV3nbfjR38AETdjdHADX
Bt5L8IofIJes3M0UhUfdNEuoMt+JrgzeP/ogscbGMBBvlgCNZYEtr8YWT3TZqVuR
Hf4L1+IXKNMc2UNBLYLonoD4dPQ0IoZ/aokXyUZQ8+kAPSHW4X+WVmVYlh1Zad5t
Fr9DtOxM3iXY5GMtX8YfsmX7YeYH8ksM2kudV5AaM+slhqbtexR8ShwB8tFrIc7u
Oa2ww0a56hUDdsntaAlXPIJbDViOz1pkr0rfva9+t96a7DDW0U/jcA5T+NxIMDYW
4szoAjc6bMdjI5usudxpLzzrujdCBB12amMCwgjFuJkbnGbr811L+GkmJdho/Owz
n0HRxuCoDBoFZ6HqyPk/EtJ5/Rf02Kmc6VbV2vpPyQ9D3hJTm1ttRaaOSbjmdPwT
jwBSLq2KAR1atE1ifOUAINcWuwmBnolHNibCFKrTghDW/ptsNbmEbpCdzNj1K/mI
j7dPZPcQ8PuqjNktPwmWFpMGcekgo+VBdkhs0gdyMoy4HILSpc7sIwfLILPU9g0Z
NxnSC97eMc+RtHiLGARo8QI0drcJeGrKAbEb8iaPvVeWwc4riPyyO+6owDKSlYXA
AwZivT9drIli3VD6zE5o5Su/sfmhafUe3fsPPSKFdR9mnnRy+HgrgPN+vcscQSqQ
m4/xlAr+AuqzaxbbG4kG+AyT3vADRPNX3Q2SGXMM9XnS20x0YrXh7nxDESWA2sDR
RWF1w1HqrZtzVZhLSDS7LnDLptiM16dY1soio7wynjfmKs+Gf+zcPe0oqJBPz2DX
M+Z2EJd368cs+DzB1Y+zOrupSMGyBrN1mC5Pc+7UfHNT+Z+xw6ypNfx7nChLEjzr
RGvAGC8SokD3jyPjOBy7/9ajEzAVuwLMSrAq5sG0mkopgiy6Z8ajfDYI/oG6qRNG
q8Wx2vTIsvetDI7m0slQ5Kcv0qEOD86Lj/A5bb5Y6OMf8ZTAsYaF6e1pY7lwwho6
Gb1DWwvCZcayjOYeI0u+LwpP/jxzMSXCQxww8naoz/qd+JRyUjxKe3OTakSWlF9A
mfg92x7j0HL6L7KqelTARJMeyVl56K+8JTp3pl0e2+AQTutf947y/fYEyJLL8kjA
mzgOzkC63U6ey87bIH8Cj3Pq/SYyWZ1/M4QUVD7MSyl4Cf3ydxF0K7GJluZ4KNtW
AIoV9JeZRp5JC2rav7r0tyA+1h7WNfYfjPBwdYHyRHjGNZMQx+pONWSIsU1/qcS+
2XXsEeFsXcWO8BsAc+CN8qlczzR1cmJdQXwS3+Mdv7HE4fBM2zPhTnJe9lqBu7ys
mNkPJd1icx8qbxwyM3iOJ5OVnE45//vPkdRT5J0bPWm6U3cBNU015CcpgLt6CM9U
6Tv2jF5q6EC3TugPAWwuUA+y9JMU/cInhHUp36Dy85fGImzd8/mvQcGrWDQr80tY
7D9/cSia62vCpo/JdVQkCLCrD9dSNTwQoYptbm9JLGU3emOs13jfEzsQm9CdgmLY
vp9Fs9JbCtSKCGTRXIkDV9VurLFho4H+q+bb5ps+grDEWK+MUXC2ePIslK61puYq
cMmlxOOfUwkHPjlJPZa+fm9xFWl2O4LZ3f6/HKiKvtZ3ZWeMxtpzPVagnGH18J9G
SujlvGbl+EA9i/Y1PUwP3kaWooJMMZpPOcCAq1/VHga5VK7VpvtJmjtd/N1Qy64E
2lCo/jQ1a1s5u0Ef5w6U19uAUGMOc4Rqhtn0HQd1VNlk7p3spPUZZq0wrjkpBb78
PG5d6dxLe4oEMqZ7SUD2iSxtT++kjAX6zK0ae7q0rb7HapHmOsQcyC4a7gtYWRZr
BgDENY41ZyjM19vMs5m6Sazr110yo7scwSa4/B2fGr5PzUhzGkXxv1LcMj8zc/fS
0NV4nKTY2Wk7GzjBNU3dDHWazrUGR3fys/+CF+coPUWnAVpSPPPzPwvSU3G7px3d
nGAsyqxRK/gZhKytJHTQqINIEU6WY2nU0i375L9wZZC9ohU9T6mPyChRy0jd3/j1
QpQUHda2Aec6RsT4cQ8+BH5SF2bnJ1A372cSyNQ73G9WfqvyMagNFlsEcp/RjWub
InMVFE8EnMOILREF3RCwjU1wiC0Kih3w5DtpYaazIC2CjoGCCjne+P4sHilUHDDX
fQs0KntK+oowOTdiqKN5eP/tWh1QWHrjxMDIFGz5J9k/gvZGeVgxjYn1GAWTGWLr
hXvkEKWSbKbBts7Djk2VxseysJOfFfhAXmyYD9JcTbKpBgI7sOn1abZ33N3+g82P
1ga3CbrC+aEzIN0RE6Ja3awNead8CvGZEVN5svirv7FM6HK6kOWrlUh0QhUxIPE8
AJs09CESdxvz4i1h7/Qvp+0fL/RBFAAElB7XCuUSiCggBYm63AShuiame5eS/775
XbFfrpEQYeMrS72TdUk0kJ1l8Yqoo8J7xVAEhknxWkqk9+GrhntnGW9LtsP3TLQT
96Igv2sULbTqOfKfkjhO8hfW/gJXEHnhOunNGIVw2Nfuy6Xef11nV0Z9WAXPQDMO
U6WF6wh4GKLYsrj1at5akk7SgNcHElY0DHtONpyoI8SYT9iN1B21xHQLxsei4bg9
rJxN1Irf04gjsKrVvLRbTmXvPigPGLB8BM1IdE7dU+uMONWeBVLGDizyfC5A83mo
HLACHtUOLldBKaNccGNUvQHu3GI4dAj7dHda7fmvFT966Ht6yksL85ZyWmldBBLo
G42R2NdXRxbXdsbYpqHHr9H9dCMkI32d+vp47krprVGgWhyYAdQApMBscyrsnZJ7
wTGOddEoGMZeKk4ScE/rlzqXJOVYQLy/KVsi8x+bulaPjQsUg5iRi8OXUfi3j1Lo
d4x4CixERng9UFng0zH9EJSMrZFBi3cfUVRTpreagARL58U/3fLaRcTeUPa28BkW
tBZewdJBqRF+11QOc4iVQrdUfHRWlutbKIyLnBs0tYVaOhOEwsxSLw4ZqAkWXtez
cbuTTmN+RR25b2/X2DCpTDtSf4n3oO9bfSu3mJl0N9jPfhAeNlTysObM+1Pj2azx
Sett/ksfF0v4nQ+ak3xNfiXPqbwcO8XgpgCaFaUeGJUOFDiNpgMn2Rmd6y9yE8mg
9u8r3X36v0vXemInrWtzTHzowULAI1U4La45IW4UZCrSuscxxp+AvRg0lONzfuET
SzV96WsRgO5m05uCkd5HyShkMbrc7sjEeZ5R18w6gvdk+twxPi4KyGGD9zRz+V1Q
USNpU8jAS9aXvnknR5Gv07XRfxOcjmO9cyh9I6jHs/gHdooOxzCoWLeHrScr6kuc
E3nbQJ5zfTOwZIWljwETAEEBRajEEq2yG8KRb3uCbyoEpCFeBJKPDCU44GuTzVUq
FRg60ChCuErrXymZW5TY0zS1ZSymWv7vvLk6+S/Fils8ejfP2HXPnHsoTyaiw8Z5
QtPRHBoQ3dJduIumcZVCd62ZomowW/TqxqA+xII1GTUEd/OEsPW4QKlYBXK+0IRP
Jft7D8PWik5wasexAtPTSe5qNaNiykL3P6QXV0GJq+VCTndFITQKoS2UymVrUhUD
NPJL+EdtHrIDMVGCarHuShtcK56zSEW1NcrGtPQjg3or8ATlUH2odjEjKeI5xCEa
AYh537F7B7RNr6t8RVILqOAIVHxI06nAf4DPix3ueUM+HfbIxJHEED6qaYHKwsc4
0xx4Onj4bfaYReQxsv/MuIfc6XZZfm4+Pt8dTml50su/dgSTSKjukZL95QBdE2b4
yUCjwszAML8dL5Lc4fn5ZokJHlHXWePp1dOyX6QpdmVtOfdCLXwTfX4VNJ4AQsZR
+4fEB+R+Mi+jKFcwrubNZL+SIxxVj4TASSM3MvbqTAsT/7HahUWVEUIq2YzkbGrp
ETg12hD8gBi4mXNcbfv0j6q5xTA5H94D7rJTVQ28yKEnywkliYpauxCZuqBE3zle
UOykUDdrKKd+7e9R5KWb2Koqn0U8MS3nZ1MPDmBbrVmFIT5ShMR/MA+AK3b/ycFw
CdUY0Zyg5AwSkIFmHw65TMb9Ca1evEitQHX72drE4py9eca6xSGMdChNWtMCmUjl
kzN+Y8Q7AGvGmTN3B7UEjGd1S0cHBg2lvzrHyTHgwFVS0FomkVVpn0n0bllApFkS
g2fmKmqd04WDA+XrjxACKnG1jXYYG1bbRFf64QavVq5UqVVzoQO/H93BcNWMCkm7
qkXNx5DPMn9oCVoU9Y/WVHZmrIxIPkk4nx3BgWy8/t0gftpIX7TDCD9eNefrfbkr
P+mkqGm6MiA2QGuIGnPDQBr5PukEr7R/dkOA+75baCr8rhPLj+5Ggv5mI3auVorW
VkUveA26kx5NXX3JrfovFiMiUWh4j8v9lL455+DiXC2eoS7dtHij0j1xJlH4DBlr
oIbDXadrkxglibePp0JNd1Pm9wpvn3WorB1vzlQJ957we9QdUH2lcVSFegh0EAoE
BtHPM0IYcO+91yQDYziaorCIjWAMu1OhqRcCwKUeMn81DTXLP88RRMraoHnfaJEx
stkIvlZKnwdVQZe5fBUveE4uRb1n09N1+/Je+fJz0IaoHRTb0cwsQ+sCboC4cw5U
QplbpiJWwyqS05w1jN4VVN7J9t1MS0dNiqcO5JWgaHiOZN5pS8c+4BO+a6j9hf2K
ir3G4CZaa1UtMDL8z3lAX0l0QBNmYJa0nlywKt5HS+aiW2A2n72LtYmDZ91IStSs
H0JR25nFAK4g4K8Bwza9sJyxX+h2seBZdVGfUzPnxpajDL/gY7qdn1WGqaudpDuM
bCzq/dOSWavx3+ZlTlMvMBR0RR1wGpRt86hNgIoSDKUZMzu4mvjQDuZk8N9PTXmQ
La1g30M5JnzV0FaedC3NgKOk4Y4CwHRsAbiOhNsCdquAKlzkNoSLG+aWQeaEjOxI
K2m8zfVcSquTXRiayL5/LlGCKrJs1CUgviOx8EJfJvPgm5z8AY/P4BL/nnhpOAyB
qrDIWiyoZO5daxOH6WYifWl70cHoIJUx8JvVhI80vcv5ZS6+feJ9OxsUQAwISigt
D1z4yyN7N0zx9bVNLiIJAwVtAfqViOjZ4il/KcvsH3/Cux8aS+eXJMwk9X42+qoR
7//koFcodJXy95XS22j1uP762Y2pmNVKQzOQ/s9YqOhiXyg4ClyuU7UdCGw82qeG
PKbqiLvE3u/Dar26e+Tc14JMhCRyjXHYRoBuMKtUBZBf4VAQ5EZXoy8183qMJqNV
9hzSqHOhfmQ4NEg+ToDGB7G5kquHnoCKIJlXtdMx/f9mPOBfIOM1haR9GafHNcCg
fKYqVJr/hbwU+RJAWVKjODxVJc1maJor8Cst6Ze3Ym8SoWOZeHZHcaFh7L3EQMjI
mplFi65oV0zwKtuuUopNaojMuvVym+aa1CR5AlEqmlzcWcDkZItkY8IotDgGgAG3
/WsHHt61gXfgqOlpiJgkEr7bnNDVtKAZVgq9/YLIXk2oJLmzCOzgCWyD3rMJGpME
I2Lq2mB1gsMMr6RckLFr3Hlfl0WYGp84cvgToIdQkQL98+UXXU/3sArurTjkHlEp
dbCLeP+tPPreR/0kdsoT/d+KHGTBMXUri5EtL0osSvbB7fyuGPv8XY4qtPb2Ckfa
oKr1QqRFB+t/GYjsKuYlgxFKYYYah9dInQr288kPQAGTyY41js7tF2vM7NNKmMZc
BRwAU3Yf2xMw96GRonnXWJQG+Oidxznq91lt86oxXA3LT5dzIgC9j6MoDP0YeJaV
2rdzqMSfcYIl9XvanEO9L6CoilVcYP9L+p+6mAYubf+UQc+quF55wNVdDQ8/1Pcr
1ICH4kAw/M+GR8eQRYig0Uy6QlPmX7JI2Ztr8N//IdBjnyfKnkmdZlV2FgVONGh1
aaPewigW8poCtRsvoc5a9Qzno/RDPlTnsnS1J06JGqyaO690q8CQz1wK8mQmsDnJ
Ej6T6eX4G14sOVvavkb5lxa73nS9KkJ8oNDCDXnt2f4zb4ygncNq+CdjTbEPzx9y
O1GrMdd9QKL+zK/ztBjYf+hxpNnG0HypNCzW0K2FhhP2d71KNVG/6GMMS14TxOND
rKIizEr8OAa/g2hsfWvPz3QCwlXu3+7zzaBGuj6bqbznORjvmBYdoYvbom7m3N5K
KyXnuolStv60FpxZ+4ZFdBaAZF5F6ZhxvQorLwxrPBDimUhJJQyKo9qYFJqEVu0w
nOpCi873E62yEJHaxFgG28yEMnjcA+9l51NmEvbk9N4q7LjRnKpoN/2Sop/bZVZ1
ZvBbHyAqJZqasZiSHbvb2gMNVxYWjQc7quFeRuyqdN1cPjYV//FY31yRf7Y/pf6Y
JcusYg2o0tv4VazdbN1tvIkKpf6XCUJWwhYkexQwApbERAErMD1PvE0kmfoMKzZ0
fCNmUsLRIfUFGVY2BjuLnJvb96kHEuFMdBuqa9U5JxktzqW2zBAZdr347OO3RD3O
YhrrazeUl4p64Pbe1boF4QnUj9k1SCFQ4TCeGBFmOO2aUEGehLBw1KnKSCmFsQFA
6nH3SMPONcLX39NQ6fkHsIoJosBA6JPS2Nco7Gw56YYfqEyIWoHDO1qD0fg53XbO
7iuxXD5e1MTvJPHAoRIeXJOkZjjhy6jZ9qhpGPA/aGaXlQ+g/TWVSd9SJH2SMzBK
2dwpwStCxDZdf3BzJkKbx+dDubgEFrghj28d85JvWwAK7UWuLAB6Mcfs4mKIR31t
N8YHlXg1aiIaX2o41ccAp7MO5OpkP1X38248RumpItGtyJEqXUHzGYq3n5e8cJTN
e/AJ1jXkiR3vOM+fIRafLiDRLUM93v9RlIZ3tsXQZShopJXhsfEhVGlLkA7BH/tU
eJXjnOjdJthFLPpxvhJJNyGykqNoTHiX6KhEOfyGiNug0/slJh9iz8qpLZcBAm/6
Oix3OxuG1cVQMwYPlUrwiRg1TF+Rbsd7YhvVzUgUimDR2RwOtZ1SQmjVvqvdRJ3C
AQhbyvmZ4KPnWm3a0D8kvYM+loNR3CPZ+6c5+sQ4ErR+OOoeqF7Ld8S0CwENs1m0
Ou/+EfoJaaof5Fc775HQ372Ma/CV++ugOzZPUBHBONk6JT8GYn3uZlIabUCDwovk
nXQemvx/FSqDJ0YAsZ6+c3TozOevrADzRNkWp/oMwg16O5LQxVsMcO2QTWD4Tywg
8UBOTI1UiTK/csoV7g3AS+ekqd1oNv7IV17oPNgKXJOpbYiPVjT4b7puLRR9i6VZ
MD58g2pfEk17N9B/bZbe5jWHnRURK4zRBh7R3xDoeBg04ggQQiKLlVF+/WXi+z6O
9p0z3UFRq6ySGP2OAbZif7rHQ146iVYbK+/BVJZRyAYKIsb7QoGZHPm0GfCzJgx5
w4976bOFoviB+5I+yDHf59XqsiiDE4DYajn9OlFYZtIkwB03/3PXYop6Oxfttpr/
o3zB0EaFcrwRi0VmxD8jB34Dhkagp/c0K/Ln2bSDMuC78nuz7EqfYjz+LdGvmxnO
O6R1fkLETUc0vvzNUFkddISicrIU3gkfAlInBg8K/AHw7lYkcbolpDWfkKHuL+uC
lDzK+RLELjggC5XileMsN7dgykZXY8Vq7SBnGEoyfbk7WaMzmBaFxdgrYkuC70gf
1Sd9YSyaL7Ah/ES0kC9HZtDgL6hhMR5WznNoIPe6rcMOGtaXSiCQDNvB2dbk2+qC
KtEUbKVv5Perq1uXRCtQD4QVGBw4IXp2eAOv7484wLDltStZt5jym+6ghInbgQ+v
vM2mW/cpk1ltueSv7HCwtJtYWWZcx21pE+8oy+gtArCWrkD+YhrmTd/jWe52g8Ax
0UG3rcyNH2dq0MMhmZRbSlDpOrBkP8kXbJNVNzzRNd3vuL8Wq9EBpyIlhFVXAYAF
njkN6G5Pbi0fLgV2reIOmayz22u1sEOR1F3FNQQ6JV9otRlhDlVpsKZoYOmc4oCC
rJht6tH3jFdllnGYK6dFHr+64bsEWl/YcBaIga3yvCP7aFcS5x/R6qYaOutgJQc5
US/Aryznk2+D/EMyF9QoazEJ9Y3etiRjmj6bl8Uw/5GEau1oIwQ5LRqINapSblop
ogDrYCPtVRO6VHbr++arGISKX9Gh0MO7Yre5v9HtERlkNAR98HUKdG7BQoPsCh2G
gi/ddPr8AlxBmYRUlbeJdoDzUxeLx7ZHX8QS85a1g9fSq1JXwzJdfIKqq+z+ujHm
rHHTRO/RY+3Ak2Nm5HW5rTKLJvvzphFNJGgxQHOk4GfcK67yogIviq1imqe/hIax
01fG7Zod3sMMbGkBn4LJnoBXmj3x9ENfU4rSNYvb/LXAHouJgGEIIz8OAALgSyQS
Fkg2sa2by83qmdFSYMRJsVI4pHUzQIlxzFdLbcxdh1iUFDJD4poWosYaBRjMCi9O
eImTcG2HgtmwMiXCMSison7E0oSo4mPp0J1BZ7StAAP3Hcp7MYKqDqIFnjXqBK1O
QUvUOdvrjGoF72d1cQiOWIYwWbpzS6RWIwZLbKzbLQIf2TnP2HYYzwo7w1FORMA1
HHOsWGMyH018ELbLZCNm7ljzLWFgFMGgAf3vjkKQxjwvuQv8oRpLQ0Ymx8hhOT40
BbEJlQam2RqxEqHYMcfgbqQ//ACmgC+kR8M3fhC8bGNrGIA+boS/Bqaew8EKY6qb
ZnTGgI3XvORdOZn6x5aiHk/GN6CehsLbINe+j2L5cufpDXJr9NsE2CjcHOKru9kw
mYAx7g0jTLIwxaWrhREtK8EXtx+2MZeJUg5xPBAHou5q/QhjZq4demUQbZ+4ZJqa
AcJ+tQCTBeD/ZQ7N/m99qpodxvbzAfnjQVggInhsJXJ512LSxcC36MYHJ+Fe60NP
hQ5HH6K4wPMWKqx72SUJgGPpHbFLp1h3N15Nqa24Ib95np47y8jjEDTmAoJIdVwN
ciAoGsqMrmT3LKlVhC3sBSmGs9iPfEdBa5pbD3Zr19uZrzC+QWA2vA3zK+AkkpvC
BSbQzyalnDjwWk2jBc4HG/I7AowdLgyVZgv0KMIlfMDP0Xm2YWvGiBGfeaDznqwC
W0vTmhwMQZYYKDRSxTxv7ltRHHnJ0UivMbBTg3TpyyATDB5rNN7vZBYeF/dLiOcS
iETs2I6XQtpCgbTuYKU9BlpFKTnwvb/+8bUTI3fy/cO1s8GMDXyD6q0Kyd6JgRHI
TtFfZXEojKgHe6x2LuvXaamvcqnmbSjzRuC6tjHtni9ZNcLf4P1L3QvY+mrWYXko
sAqHtHBfeuKZoFxp/2LgQ1bqK1wWK5iCH688TdeyIsfSPQct2dD2gXrhENRiHaCy
Eq3Ru3oW+an0PvOr5FyGTApkfGOkBkOwdWBEx/4Kni09XSpxrbmM0HlW4RMXkBNP
pO3qbR2YXQvzdIa+3n+6qNqDdA4B06cmVX7BPtjHFO00/Bl8vxEAe5IpS+9sUuTG
a06C9TP+AKfRPJ2KKMOnfW3XvbPp8ULJ0D8KFHHMoAaFY2PB2tfJwHPqcQNbWud2
qKncXoXTKmOp/EDtP/0j2yjTQveNkQTFg03OV+bHHdb5gjX0JpflmVXKNJaev2Ky
GdoXt3FWPJxbGepfaT/QrytPKqgU3lPQLj9ezvXkTs3j205P0gwNEmJTo4zQUd7b
F/z5O+jC7J1tx41+u8FrbXUo98x4mxO95stPJTYr3FhiLuKGcVgE5r5FJ0KKlaAY
PLdbYO8h0Uwx6PzaWsw2eJJFr8aYtspPW4mkJl2vgzFIiTvhnc60na6YmJlcRkZE
gdycLqr0DcCUHB7Hor74IwfmB4bAbYsIBRfyzk3AuW081SKz7IEw09NV6dn2SePT
naftbipwe3Q9Bsm7bW3I0ER3Jz99gOJWW1oQ8+xtYwqT2npK+HfpbYSkzQ43HgHT
3fskq9pMNCcai6Z/Cj4FWFZD+v9qWhRJ+7FCro6c81cXkryzNc4M8agCbj9S+KWw
g54d6t6Bq6L5BWf3QwsBurlE7StyI2xs/TMIF+EdNvLPGkWjtuVDarcmbXK1Cmuk
VRhTpBt8Ayeb6qvLYqVi8DNC5ilR9sL7Dx7Yyrd/JoGyNF7dJacJ+D7PBhyo0ZNE
4eMt5Z+vQEr72dh/SlOk1JsjsBz4xi7rY54OD9Xs9OfOCT8bckxhJ72EZDtjVmSQ
VyDzd1xDd1dCM7Ykv5gPOWWWLCuwIf4SSzaWDp2LB+gVnQkc+VhjDjldvCQAh0A0
KpmCsgaUX4abDTv1uVoJwdqmUDvrGx9V/jVskMqED0IydkNT7WbVeMR6hAJwzUET
lwvtoHHdQhvrVs0ftJ/wcWBVpziagPrgPPh8T6mIxDqSJBElIa28gM2XPzyyF69y
XoaZSq2lk0kCsP42EPw9+2qH2YfSejTHCf7CUnu2yU1zmr01nl57cLxMg5vzIuQf
vXjOXxkVWLuAbD35kVHQbquiq0WuZhSTLaChgbqDlGZ45Bv8ngKleQnQtkJaQk8h
Lg1LD/O6yzmEq8f/RrX8nV98A+AJYRmL6xCQEWDNvfK7yVkuWxXV977vkzY0v9+V
B0tHPYDN/bwQhK3bhA/YdHcSVt2+BPluat6/ubVJtl3g9kRoIclzTxwo3co4rbt3
ccx6GQb/BMXMqmMEBbvl59v6I0oeQe26tkJHtopH4EP0FxNWGhdo8jrtJwLh4caN
whOI8fwtcnmdDJxfEQHagYbMVsl/hkFb9gDuBNe3L+mJ4+FKDYBnR3ix7igAj7fs
o41rzMRs0/v9yRacizYRBO8S2DvvIAAisxnyAvcEliPh7y46JW+ytrACShmanldB
zx1wWAFhAHmsO0OU0NsHEXyAN3dCw86gB0lPaV4xnxo9hgnYBtQf+98s3eX3dJus
LeMttFEsnOowYRjQI63gofapGdsMGYyTUrsTwu+u/0ciucIJ4/jgK0gXoNqiiQuM
E4YTRpYteQwvGg/n/sUA/FYTkMMwvq9aL550LhfbvnLU0TznV8W7NXF8umZtxf0O
r3+P8gKeIIXj9sFs6r5RCkl637ikM3GRDVtamNffrAcZ4joGxdSNJvqAJdw7FJfr
KoTm7/bmvhzK98cuQM2rrhHZydxzONxzaqJsRAwOAhC506iIVa0xwfTBcf/hz4pk
qqdzI+1lK32tICKyoW/oK6HMRpsv1masSf78rdQ5+7VhHXQa+cgMzvKdwt/IWTWR
lo0PdOaWoeU/bIV7Ca4YQ5wXUFaYIRhbnxteVeAIwB3Zi+aZYP1vnJy6BTtotqkH
tDd6HvTKker2zMiilhL43myjcpQB1g3fCn5jLokX+SbWjnKGGg/gMzTQWwAJ3ezd
WoPtKufPbp+iPYEgjD8H+5lAXSUaTBYA2g6ODyGM/oDNEMHHxlabdxXBE9v7oWAJ
0AWfCUHqMBnyhc7m80MSVP/t0E9g6abFid0NuPsrTSQkt/J2j6HEjMxBlE+fhUJl
K1pDgb5krBUhXMyj6XRKxmYqcJayJAeExxoiakV+X3gR8e9XaLz4XvSUZXXaiZFo
HhJ+lq4sgqj8+w9DbQUynkt+iBEIB13QG7Qqc/W8nfOg8DerN1TSmSGEpO6Vj3Pq
Hpd+eG3cMwTK4QwlTM9EjPpQTajg0rVX0AZISthRjbD4w3/meStn33p6WfqrECYl
BR12+BUG432M7R8T1nUBI7+dOgn03mXGFwTT+B2JM00Kk8+q9KNrJqdzZxlgTFWa
MOaNV2L1kNUKMdzXAccOSNMoF8tFOcur9aA2QYdyy2CjaombcKlfIs1UFKV0W6XO
IgLoa2gjgB2dQ1Ak70XHubvxn5OZYtVTDZmMW/XnVqpFfVoLFlM1+EFoU917+Isc
2koKJMiUByFgykSL/zBcU+N3m6ygUoIxM7bzrlXGJSH14x/y/EJRk2+OjBG4yVqk
tRZLMaUp8aegij42TLyclQsgVAjGiCbYzjW6jh+eNv7Euvafs/04B9W5IkZ+rBa9
2sI+DeSwEa+Csz2EyWOeoRNw+5KTeoQd0YwET7lvAaS4X4hgLsISFXNoU0U8ZOrU
7pzcT04Zr8KD11I9UDt4ppRC2ZS8NISePPg1J9T2WcWAGSa98aBXgo4O9dSL2REt
nV2QCNnMUvNkA926Sxmeg7XbyDKUqlOK0f/PhqQmURZFnbLmDGaefa+sfO6P8amC
7i1zrZWp/KCw6P0G5ScdTpz0Sm5KHcHRSIlkaaZA+yNoOLQRGyrNs13aDEQ1CnqC
mB+8R361clZSW1d0QYn872My6shPpAe17BRAen7GECDFeivmmvd0XAmS9sBzyctR
oBiBUcT0kRmnirFvuO2KfJxOl83MNC8qjKxPluVNUoyRW9wlB6jkiogHRQIPiLJQ
uKoxeFX9K6ST7FzPo31NxFgk2+e6mxdPrw3ljPd6vsfg+buMpNKksKsIEwvudOXW
Alopt5U1/0sJNE+Wt726zREbRRtIbEJL4Nt5hcxggwyUr19HicaGngh8H4Fl7snr
+bkN+9OcOWKT6vML7oef5fynsyFZsq9lH2N0dEEVjPEyPu3LTXAVT3GxZxCt848A
ag/uZoS9tc9zW2F5cTYK/Oh4pqK732ygGhT6DUmoCKPQkpavAth8VA2t75bif4qO
ogaT0MdPLrIkeXWlVExLOR8Zcj8oR4/U9ahMRJmXC/qs5e97NlDsiB4rh7E/o1RJ
66F5YKd+C9YIpHOS1R2oOrfeXJ/OOGTy8ihjgT432EaZ/NDV57A3AgedYeWmoCs1
a6hvL8iQ7DlhNTaYoUEOOvIm3hcwtP3l8Eq/igIRTYKbFSQdI/huNZdfUcUqZXHY
jOneMxc2yB9QqR+0EZ8/nWzSnvH0JOR9f+KLB0Mvm/mQwhve30+qLuLX8gejdADf
TztI0k5+RW3fZadK5oPEcOVKywhksj3kcOjYIaoYDqeM2CUIgl5dyN/FUCqa83XH
02bu7OEmsglbzaCq2cwuf03midSk8eBhKbf8ppBR3/oJ/eH1xWIFkyDRngL2nuMI
It4ND/TrZ1G6YtX3FhoXftj4tCRU4tFB6aFSSK3SYmF6mITeLJ5q4/CFDsSSIMb6
4CuNjAEJ6CfwY3xPRcFRRwODTJ79aSPpSGhgV34d0ud85Ln0tVUiwNwC18pZprbQ
7Y8RkVRrHeI2eIfToaYoT82W4dhg8brK9xAICxRIwRanq1SiWA9Uzpwr8XWaTLYw
n2IYxfUskUfvdOWbtUmrQZ4TugDhwRKdkEAAajYtmU6WKJkEredg8m53S/q0DWLR
d6RullrC1tof+I0s6ZMkeNNWOoyeFsx9hm49PE193iMV7IsDEOw2S+JvUMrkAuN2
hWxQDMCVicnEGzxROVubg/NiXWTTCHcLyc/Da6EeGuyr6KVh2oAfDKRE2Kk7PSr6
0YY2wivpdX/7SW45QbW2a6+0hwPbwGmrG0t9qauHqInLsbAHZO8CCEF3I4pLnHqt
9aZ1LcYfI+bTF6bk8lkEkbmESUtyqb/E76/Kt4+BYGARYteKwsghnT854TC5iUdU
DF4iaGxBanRWAt7eHrgUK1JAA677iE9qySSifhnN/U6c8U1CqO1Y1JbRLZA9XmN3
f+QcsqEllfl4TSCn25Qa7qdRJIJF2cfP1OqOb6UdBXMZAWtjYcY2l9w2Lo3Es6iy
C1hPCGAg6NUZuN5uB9OfTeW1iA+Fg2PjSk29i3IrZTnQAyhyHlGLSQLRLcmy/m3X
6nyUNYsbg54GUn1N+949jH+p3KH6nHrnkskaPGJNeABsu480IlTzPMfwIJY1MqoM
P8T+ABL55oHuZSWJytvfy5CV8tEdtWfpqkTfAxqU12bFTPunXfrHOjGYpIG9ufMv
n3gJv2/aSjuEBgf9HQFTvtz7ztZYEFpEm49ABViYBT5W3QDFYwG5M2u67cpyPBMt
pXFfIN3F0rc3o6EVxip2iVynaFKwWIa3IivjIJ9pNBar/GHNVklyj+w5K2Bj+Glm
mjQGVcht5IgBydNV5WXh4aA1V13o7caX0cIN72nTnFZVXVoKaQ0Kkd/rEBk2rWKd
HtIS3ZBLr0X2DYh1KN848nFn9LvscLdnIV5a6rSN2TYB1R1Iek/QtgDywouNybGr
ng09/qPM2ZvxrIOat86x3mdi+5QniEENLE75YDpkAzYyS+1vmn0IMUPQYCWJ+ZNU
1ndrjLKuyvmSiFmGoJwoNFnMpf/etqeLU7YzQYpsrHapZKaH6E2hyCYZryO2h6TY
F2kjD6GViw2l8UDphA4jAJZh+KvEVPnTknPtXBbnIWo5yTx0He7V0zoNNC6EL31o
UKvwdzcpaFj7Rg28Vz8SLqQLl5zQ8ldo7o+tjLHdu74XPysWKSea63QDUzQQ8hYx
uEolPnqOvTvJGc5UQNffDlQTOgeoZGZBue8OlzQf9qT99JpXcYsm7Ox7oH+C41QF
+Lwv+oNCuAeo0H0OIhSXl15WinWsUJl9pHdDGcRoNxgzplMPdX9Cyw93zgcYtI+d
D7cQjnrpGI1F8+WheEQ8E3BTghsOxL0uQqd+hZXIw37eYpxjnAdOWXruWoPlWHi0
ze9I7EvlrZaIzIbxs0wMWUM5HmUReale3abyXPaEWJ8gyFF9oevF/+p3KO/Lokjq
uz3mjEOGSHJ1PePlHAkfq+dYKNrgyU1q9Hvm7mr1lV1HztraSvscUOR25ZGqmfx2
SGwTYWcHXNffILuwUsbWgKStlXPCgpfHTdskFvlVamQKd2yvtQbyhpb6/oehroNI
UKNY8TGaLl7Ys5aqW28qLSUMOofRjuddO/GT1HjP5rCiWsY2/qn1nIU2301K2vyQ
SsinlbWd5KNBv6yZq7WZz8zudE61966kyPCinTR7Ltsx483J57qHxn5QxD2g5uHV
Q/WoN6igZjx+gxTm9ShUYqy5czVpuVijEWNTR0itgXdsxR/UZD0UQ+xXurX2iHeO
foORtEbU1FDmCkLVHykQnxd5m7pt6kROerlM9XStNx2rvpTGULDLSk2BG8KnB3Pj
frsDZm5r1R46InjZ6KEyv4VNFNQmncWR9WlEaXxvvmJtVhN52e8mfEF/zE/s2Sg6
XIefSMMrAYq2IpuqugIJhIleZ9Ah7ZT4g3NqEs1wYEr4ARR3uEQh/oM0Ta5ogbWR
rBULxrmHw6k7EDc56jX6nTPLc6YyAY6jqbNeF7DMDHOj/jVuc+7iFp0PEMKF27IK
MD5HP+yzMMG6eGwB+XpKHWcEZCuSDbg1TMyc1XJDBtb3Wh8EmcFrWCPHQ215lJG1
FMfXY4X5y1mGk11WTVrGhSxhsdF6TSpfCs5q/zR+M+Ha8P3A1eucMFE1G/JemnfV
qVGyYWxcq2HT3U4PesbGz9MtWEi4l6dBoGTcguOyQFM6bULyIr7Ey/kYgYGBc95s
ahL9s8bAuSD6DnR24o3UdCvJHMdtgfVmpqBX2gajHsDMb/R0E4MGEo0Zu6Nphr9l
8uO2BPAUEfRt1eBWJvDgQ6eigqhI3qQiohaz3oxmTNXzcU1YVwsnkzbKksdiL5zk
wVeboItbPziHrEuXAFVIZd6wZHW619/ZTW4NwzcECZw8ZFlHE0J0t5fsp0Ofha4H
3QgI5NdFFwZ6VDPnWI1P4Q4EJO9vpTXZGMKg7pgegPSfW4gTSOSXYNCUd4dRzN//
JsgQ8BWjajKeJask2mCX4POm177xQKXDcAN4FMN6OWth4sgerKnaLqEGgHyIfHON
X/mMqejz2H0IVNGVsZJmmX8ibei/FQoO8TavyMtIYRRrCkxWQBiAeqekbwTF4qQV
vvpC6tnsI884WsW/HEq12vSpLuy9OykLfWQB6XK71TaJtDicppG0poCFJDcSIqEq
GlQ3ZhK/VQhPWRZP/qyr1u/xLl2n3efd5GES6SHNtPLjpSG8zyJBW2d0NEke5SpG
JlNYlAVtn85b3LwQW7f8z7Q9MyZMDlRk15btQSODkUfBXTBRAD01VfC2AVyo/uEY
rdE6MYDiuGaJlWqOFNpvlKCpeUvtLX1vvdeWRg0IeuM7uG1DkLfdxrplXAmy8tub
zYXTGBSFLZUBgUejhI80R+ze1ndm2qgzFJtUFtpGqRpCABWMWKARKhmnQetHMadF
WR0LhoXGekPJMOI9Gv1oNIAF22q9MTNP+NxDJeeDd97NLdiGGosR8WEhnFv+nKIR
0wsecJCEckiXnf0H0WpKct3LdYYT54U/IFNlLBXpQ+fblfIGpX5QWLssDN+Y0pE5
KRQ6JP4zJnv1mxigPy1ccakq/MfvD1nOi834ag3qLtmmt70jDFR3yvS8cPS/+8+p
rXdeYDfXFsoIub5xVFZZmuvEAnLhAxC6W8x4PZrrnMWXjFw1kDBg4Oi5qMcRvM21
+sBgp/Z5tB+fcKh96cDNC19BKwkcSL/gsqsnNCHSKSq6z0EqfV3xYeOou/Td09q8
zCZ/h20+isTCUaqbq+DGCx5MSzXAGaLcZyonqM4Uc+lDfCe/6ccYpOe/FO8fy35P
Hzxhntm+xLa0g9LfGItur2pAUPHZ35iB6SXOvnsJ5C6I1jf7JsM2CbplfYregGsA
mnGOGFk7Xuk/f0nW31AHR/eJGGkcaMkqGPsk1ChfJIr6lEJvLsGyKUQ8SxcewW20
0FBPTEggPrpC8ROMh1LRCvqpHOWGVOrZmah4tianp/GMXSvsnyXTljzPeWtl9I0n
+rzx62aM9qqhgSNXtUj/NNIoMKGSa8o7q5wwWNsUaiTmprWtBuwXWblK2ikqFcLE
TzEx0qafJWrTKcZbvFp5rzcg+SZBp6X9yAKvqkYCVj3J+LpIsEdnl0mSjzndnwYe
XS+lfHMRlvssJQmOuzBRKYplrnH4tcLS9PGI5X8G1CWzRVQHNesDhINuXI6C8QeL
4Wn430Qxap+bEREluiU5Wm/s636sa9bGQX5ojwiXA0Ie0upHZk2IajPtfZcFCb91
n18WSJH059oq6X/PAQ5B7ZTMu0j6u9LTtyDd2Kyg+5urGlH3GF0mHDxoblovIFei
5pjxJkiSCqXtf9O3RyUuJ9uoRQUtf/PFPRDoB7ZKsOg70znkLzlbkZCUTDO4kLxg
sQSlw5nNir1dE2ErRUflrLIkA0/dotrAhPNPjJBgd7cPJheYE7L752nHaXKD2ECV
paMHAahCWI/vJY9vRRMwpnZKd9vgyJGkemJi3nAOAJOnuoXlFxNBiYo7BF7Epm5i
ZQazHLgJZtfJMMype9lY/QbtpEGaPyQuP6xTuAyK/ZmGDwSDBDNnBiYrP4EzBLzx
6EzO8Stc4OhA6/K2h6Eo2NYhXrHeCyr2PzN07fDc05L/ZnXL4OkEOR2Rm+KB86Sk
+kKIsoJugKIvenbQREyLbsfxos7LuXLHzZM1oj1vDzTNHMcGHeYNOR+ZbcX2P6dQ
To7z4grLXHcCLaVboEO2qYoHYDI0ISwSUJulnhyu6roT8pZFhGT52Brq915euUpP
aVgnFMaciWfZp1/idJuu+pTiBFDBVvL4rTMfKcp3VrmulWz5H88W3sA1qqiJ8qOA
+ColwqBEPKF5o55425gW/CNLZmx02rRkmV4NKwEyArkJs0mQFttmDt3QBl0Ybe8U
DOqy2Hmz1FEV4aqDe67Th2Hca9Cz/Z3u04tdorE6ghCdpsJsTRx3L+NdX1uAi5AO
wzUwNSGhiBbEiQFs8xRP3NsLI6kUtVB+ORe374eqrNij8QUZKOyy1/0WbrPtf639
pBJlClNtYVKgDbT6faXjLV5m3ZaB+/ytKNXjeGUydoNs0kkOrKj9QIS//m43H3gy
xrz2C1doF35iHmhdAjsx1R50ydavSIEed3G6/SlOhaq83s9TlonVpf2TRI15xCjX
Po6Xjn0YVu/FU03SJ4XNJaqeXdxaFOHcbCliH9yrmvbjM9NS2CTgTJLd1nQA9BG0
YwKkaBSaVvnHCwHSxap1gyHjhFnV1jDZ7kEPmRHrp7TSYy+ctziiSI3NnSQZ65ac
B1ruhPYGHQEfxDH1VjDXVhInm1Aw2o2hXhs8AmrDu5GyT1dQDRCaz/s1T5829shJ
ttiqY6CpQ6cENW7fBASanp1uzbCOeEQyzV3wc4zGVF0rFG+v/VOKMuMyycJAnnya
ViMwRN3EmhVJv0SIpcJ17hLglodtPlJvdZ41bM2K9w+nPbrawltwZliJG5bg0x5Z
mjiqPdNLodpgMr4TF4UZuai1U4/VkHt5duXOvDNAEdaA3yWIwjolvSGI4P3se1KC
B/anmMfaPesqswlP+RUJ6XjZvGgrKuXC6fTaXok7EUoYseGQrWJQofrAKWywjKoA
gvZP2SrcoRSMkjsxI0AZ9CLS/9JAvUZ8/sTaRvVajJp4EtNqGpxvo3BYwILraJFC
ylg8M2JAKALfe+e9akBDhnvxUVFjscd/w0sWrV4L/ycDO0c63QYlB3uFItiXp0J4
emsBFBZMClna5V4SuydFpaDPwHx8cNDtlXRzQNDEfTcATMISLwIjkKsGyuFHt6L1
EPNzc6T/5ZKRagptSRW9e3VGje3VUxJk3p5REtZQRpAVkQSp1ZAeEM15LwCLqaOl
NBYF70hBWUHigzXhAfPZ8Mq0yoVj5vGf7wQjNcEOJVpPdHZHeiSXeAR7wNkDjO+d
kC8T81cXwReJFoi4YkvGWiSt688FvTatDILRazN5/9tDKNUm47JTVLZOUEXS4MbY
f01wQ6xNBPiBKt1OEKKObP/tykHTU/aCTqhQnJ68yGjgJ1F02D1HzFwOdnmWmYL3
RKh9Jn0Ck39kc7so2401OeP2dqP5LRfYuANz4n9dGUyT1rbasDsQaiEQ3YeP0R/+
ChbwWRWHa17WUPlb8j+Zdh56c0QCsAe/cI3PdRjIuz+91Cf/s6wRmsmR62UlQoyE
LPynLYOogmwl2noAgr0zc3B9HBvfMFaLE/zhROWieACgg285SNvMt2J+zQvVEzq3
UIxtd42cvoq/8MiNL2i/VK5nDtpHIVhWRPHU31sHfuc4fGIGPZYoduvncNw3sD+i
mn66RRMIyuXX8luSEYjgIsBvZUEu68n4dokEMLp/XCpNSkWOv5icDd+9jc5FwqoA
a/FKoXlWG8bq5U+ZKfhZZOEb9r+eDzOVubMMz41vSmraWOf6feYrsmDVohz9zsBk
Ah81zPmrWff5SALXzxnVIfkzVWosMEmNmFKSUjJgCqG+OxabIxGA3SHC3tcXyrmc
vzCw/XqbztZzF8qHYuE0SKVqSU38Gow2nXdLHa3w37oE3P1vIUqJB1x7Mmorc+f3
+TcTLCwx6MPzu6FkZaiUIVwaDdijIBn7/YmSM0637pJn5LtXUjdB73yzp8soGzXF
9rv25Nwm6pY8MAThPpXqrGP6A2ktTR2EIUhJlI+in5aoYFRZAChHE+4eE62Vsndb
H8w9QgqM8VeOsTi1PHToAJX+lNLwHZ/MWljgkkrPq5nYIOIe5oDT+v/UnV9qriek
Hl+2Rx+R8aDlv2zIEy9Pnk5NAfP/36s4rn5rtPm3xjXN13NrBnTuhtrv9EUNNEfZ
2z346jfOnrqcR85zjylgdDd+m9eU6MiQX7PZODNKVNY7kn5t8//er0TF4KBYpSMf
ZanNVc/DOxQCZ0YVdEwpA+2jYbMw6f16I9Ybuz/ZZeeVG843PA4WPzQuU8rKcIyJ
GYxmsPMbrYKEk5/KWuXWpiFiR3B74FCjrvohGb7sSyUgymIlL6GT3uwzlrdmEoq/
5eauSiXeJP64e0BLw+0i9VlhbRcICpMrN/CCPI1YaywcL6qr+BtO9oEzI/1wGDmk
z7ICjVYfzWM7ib5wDAKZKy8BlZax3caaj81XuGmuH3BKeMntvR+oFDACJrSXi7Tx
uAM6N0YQ8i1k6oDMDD0GIsh4bDzlpVzAz7JisYZn2vVRfHM4zAI6oxLJl92ml4c+
eaahqf7gKaJmh2lw/jgVG0TzXiXDcL5hIdrm+1K8PCe7JgFWq68z8mYds4q9YUeI
N6aqvst10vd8N78tSaRVy2azreVIoSNfoWoR2PV7/4QsdIk+/Xwm/q2CypXAyeBp
mM1gzoVdu14rAezzQBuBWvvuOR3m51OYJA4h90GnobD/dVcHpDoN7lpgCDVoti+i
Nt3QdU/WsU3uqLeuwxpJkOZtvReIOiovqHX7ZHnngapzLTvWQ3yJb6QXUozOoVUs
oqnzhMg0pDAC/9s/c8AO2b7Ot9nbNIXiCM0yCYDHkO42S6ibCD2NcjqASqTDaKSE
gtqkdFYzCVg0li3y9PKhauXD3pg/2f5eumobNkTc3XN69NhyANyk6AFgxG/n81l2
1xKu/6jJl1u3DZuvUWfkV+AVnWT8qq+RkRMLViGy/nuq7ZsoZoig6oDL3GBBcglQ
iMh3yHcSJexHegKzKGM0eHp1txQRbWQqW0HwTr/7AH+B/ADZvyqWPUgzDEefv5fY
mhygm20YoRoSqAtW6/IbKaBbx1cLHu2IFU7UaUDO59fjpNKIhcQH46Q18k9xaZ+H
u3kVFeocB9ZXQ1TzzTqrrlifRdhcifzTb+c3A2qM8/eiDnc4CnZj/LQ3XrrThuY+
LahMVy3Ts4lNs2aBXg3Cno/lyT8KqqvgJRx96SOzO2YZQ1Nlh6mgUmwDVOCUTo/F
mjmgJ8+t75vXXEOEZFLcVi6zu/s3C3GdVqFHpiNbAxtHqVIbOGGRsJPAhapdLt6W
+wbyMF3Go0o+qdQ175p5q+KUHEASvEH7zHg/031cA9C2q78XeWUGyqh3B3Rm0GA2
NOEKGoo/5VW+ojULVgdCj7gCTSnaLw9+XGGogeuVDzjwwAGvR03zw8XDNs+0L84D
LZU7auxaB2WUOjKOtNGtPLUqDKeEuvAWapIhbrUryJuAP4GICROozOinvY1bdmjf
dtyTxeT3jofFHqjgU32aadSvXsYExCrk6kqNhynimLjpQKWe9ET0tJrx+lYPGFwn
M+kF0etm/IMPHqbT1twpMib3aYRQDTNxGUAZiGHcSjojHGCax2pkA/N5NWrEW9UR
Iq7rNkn1VyRNncRryPDfxogDskPTeW6u/4ib+adiV3xzNohyxfEN6v7/qdP5QO7S
4vRu2D8DpZNmEsDdicZUx0aeZ94Tb1nBJjH4rClNmR78cLzfXadiJf4Ucdp0Ardg
jU/7/p7e6YVLADkx297ZUb+FwnB34wND4lWNQ4vXqMDXKLZ0+0PMazilKlq5ItR2
04Blpgh6of3ynTGtTPXiTK4Drh4lTdta+fiOGd5JmlbayMhOeZiolCo0/vvo5TSF
l3zCRSFX8f2N23UBV8SKsncpEk2ws4UeuGhAGiIfBsoo1dsSMKFa2U1pflQbTTyB
Mq58p1BRuMGrw1JOMSttHNFfHefFuVgi5720bBPmjQtk5cvUVLaG9qSK6fXUsPM/
beYLtrsCic1IdBJWVKvWJcxUNBoOj9OZCHFcBy4xaWr4zzs299M6ghGokjPG/RVz
LY/MrBPp0zzkLsrRuvAnZpC5HsxQtECue2VsPv7t2pzBBEO5aM4tk6Zp0wvbNJyx
TTAoUCwi7Nmg+13C1pZvNUrUOG0IBQLCq4ErqcHR8mDYs4hs647XBg/9EmHu9aQm
wR4J7zrrpJ8vHO+P4Nc3YgS+J17W5Yp2vYrQyXltgSs/IjXQKR7TIF0o7io+a8fR
wiZgL4iMKJraxgynU6tSGkSftUKh+hGFPQH1vFDeWlLRS9ahli8v37cjXbvObowR
Df6y5CenETyTqDBfQF17vThspJyaHAmEq3hK6g+e9LcwqijqBYhtHXkUOMgyqowT
KlC1x98CfWsdtaHT0KH7A8mV/7co/rZS3pf+ALLINeu+nvCSqIKQ20d90hN58WyC
KE1kYvXaLVqUYw2j9F3+k10QrPJPoiZeutKdZ6nli3LnuoQEXuqMU1BoBEzmqpyD
ZBnHU3ScoOxzkgBCgOPFPbGR+yCMM98bYaZ3ffeOBZx390j8N+QNb/K+RCzklN3h
MWIbt9fMTvsiZhex9V/tEYNByeb4GmQIK2r2fusaAjqMps+knPmMdi54H6HhKviP
WTh3fLw9MUaY4ErmqD02vqjLMjHdAsvcchZyVRJA3K3nK6l18jkOG+Iq9Lis7IY5
XQNF0Sgh3bnfhqO8wfF94Q9K/fbHfVPxa6h9uM0jEu9TzC/wX6hQzjrhEfdUX5ul
uQNrXHnpdx59Z0BeXWvY5OmI5SI0oXAsEEUcY5iRWVeexmHa0s2hc/o/UIRfZZTX
Osn6q7ZIn66Rvt1RaOegcWNYTbMgb/FMo0A3N0fZ6smEoDAmjRFgmaI02WOUiE5x
BGNu0yhvssiJnJ+vejERZk82qbvY0jsnie96RX8PjhR8s/LQ2i06EkddJOKJ3DZN
NauaKJgCo+8mbHckAwbsiI8dT651ML521YU5tfSRV9kTg95XInOZfqBzOQa6kWg3
FQvpbxQ8aSKn0KEfJiRwsIPFweaa+HgOwf3mR3YBa97+fDVZWOwHqoLDnF3aOrpc
kgwKVkEnABTdBoI54vRICdzq+edqXvLZEV72tKH/M2cx+xaltBOHlPflKnfarsSQ
sPDi3nfDlhymKHxrvCwZlDCSv48xS/RMcXm6xx4OuytZdx3VqJEKie72mmpoUZkw
lNIJC6fRNwyHMYtrMSIEZVe5Y3PV2xKaHQripCxtvuJJQsYDgyqTZuZAU98aKMpe
MCk9jCe0uhf3Sc4CDh8gUIW/qWOH6+vk/KUzCuSg5LCnsXaciuATIw7LFRl34nwN
qquIbmP+/Pex1hch3mLZ6w44I6D1sDflDnehHXE8QeF23hB0oB6PHY1v9hTfgK/k
LLi0b/IGBtSBsoFa//EGjWhuT0FKA8j6iUf4LTosR0RTPfhzegrUaCszMxbFHard
MohTh+FhncF8y9mLrrNhD1i3r6cb/6les7xDUqg33u5DZwr9qhjy3Vz2y7wNI/pc
LZkk+wZBeJWCuRc/drHV7zYGZfh5RdhyTZxShHGLq7s9nFds8MCvie3aFJ7uwpb8
UkAmI9yFe3exWFRVbiyf9iafbr9c3MrGxzqP8D98AFCqIPP7jvq1eZnSMRRMrnnJ
omcaW8/jRjKqbRONJr4GrrQJwlAdPlHAlYCHJKh/PyVvf4lUSWk+QyuCCca0KowT
Lq6CIoTouHPVZF5G+tpnKtkCoapbeTe3jVg3AtYsQ7LZH8xVwW5M/LA6UjFBEHhG
wn40vnwg7G94ommSptCEdAPmgmCS/mxszAsKtbv/zZbuNbI8EeXd2XC/jkMKn7jc
SQzJkDGve5PbH0HUrUKiU+YD5mQZTR3yq9DEBWiU38rr4it71UpUu6cs64u+F0nf
Ycuo7qY7qe+AZ8rmSBBuSpzXUg1OvbAurQG1ZwWEBfk05IoXICEP1OQTLeW4b9UL
WIFAOXyy/+wsxofuS2CbC8YA5XuMFsUC/Ep6k5+gXT85gJDx1JDRW1wQyjpnJNEe
sd8sPPokx1tc/8Y7UYGTO8gPuERa1uilosbrPPgNb2czCnsMLsuqqrQxctkJT22I
iOSCsvlwm53c3B3983srHrlwXxtNnwsUMLCiAv+GzzlU1jCd671pOTjzfcDgl4m/
lsCldAzR6xvpKediU4uujnxJv0vjS2clb3OXmTd5wumnc6s3BXX3yIwlWuIvUmCz
vODG6G/y2CNRNEc9t8domXaOTVu+M1v8PtavxrA575L45MsDkkWosywgI18ReyMe
wZl09M0utlOdFUdTSorqXgjBeKnaL40+gU9NWbVbwQydfBSkXuK0CjyI7eKf6eVE
orQATFsdCsYZNIESvgcDVYPpCs33EaVw/eZPSEAueV///ENMZ0jorBNxY9dzXZwq
y4lgyiJNmsEBQdXVjxM3U3pLPiZ9ItrVlESWQ9q4/xjTaEC8Kpyx7W/jE4gJeorf
7P4qCj5YODDR35OFjz3VVz3taQV3Sg+w3HceIH2YmFsAE4+6xEAcu8RAMz4yPLqI
f1CDldj+DjdewupNv0xpvwbE4bGyDu/uYolNFdAWMgf6gbfI4M5qbXURsWwciZjF
yTNhOKMOBj8nhF3jc/oECMagVl2FUazknxjoXLPJkab54jo3pmDNkq9oOQnJbi5B
jgpxSkSVFssxFLI3aEQsYo3RYYhpeQHKznuYQghqIk3jml60Luubz9GtCyONfFN+
qa3UU8QmMDj5kBUXnxi5gzDL/n8B9scjgPZYFKbYpXVR1A7usC3j1fghQMOqdTEH
ExBR3gCQfwMQ7qPLKrA3K0Bpr0kWRhDtBZBU26EUXPBixwamC/F8OXsUSySsxP/Y
tmyQedaioYopWAD/jDoisgtw/I+NfZuTngX3xBJZpSD0kfZrSZ67e7M7+2PDx+fx
YZ/bKY9lR6AKEXQ/cgp7HezgMjnGxR9FlJfj5YPcX+t3w/vQ45c9TQ9jVGNLa0Uj
RxQV/GkloIWEhhxyBf5iCvpJD4HDbitfzRdzcNWTcxSb9f7kfjkqVfgYWCOO6kzf
Rm0UgbIbnESb3kqFDHfjvcWN1IzpcLEx2Q6bkl2WOvXt8dHYYEOzW1kxEDtlVOSR
A4eYB0FBZdaFIfTWe250duwvO9bbzbgOsU//BImH1JWVnmgVYILWqpLWqO9+T7Fz
nvhAndyjLK43LJ6jCMJdIuSeFhlfJpz1KOG/ZcQvx/3yIEnGsQKqHRS+Zo3HSw1D
M3X8Ub019EbFvWKz4SxKZbwneyjIcN6VFuRYkxNBlQv/G4UEbjaP7xtdxLc65kGT
lzMBQT6jbRoM+UPNgXQqj/25/vRQ61jc4vo73JK1huAWlLqi6X1sA/rYZctCi208
xzVYcJK74IHauKXNN6hwh2EjkY+Rr28h8bxkicCQEnh+cSchjtTruhC2pKc0u+wC
mxGeShyIb8a/HsQQDdxmxfStMKJJbkb4dx24PZH6C998HD9/8rmkeq1bextw/c3+
ciy+FTF+FcIyYD5I8emQVIdenxjAXhNnktckNyeKC9xjLRpllEHe5SEqk+7htKkW
C+laHGoQ70A2WLrZR3IgsvzxDfXAporTwu/3V7+5vudKzy7X6mJ5S8KueCnp1CQH
gn/Q99XFDELIVfhykluvd+5M0CAbcfMC6qrpDl3bixf882U0/y3ctNWA9h7uTqv5
kjvWPdXiPNTOpWEs8zCGxFstFYuu9e9h7z/IMcWRlLtZQFAbehFUfSRJQfaYdl5j
RJBEVZvWVwkt4SOb6XYxsZtVbO+DTN/ZZm8jKHI8I6n64LXdSr9FFcNM4IL7+C8R
NisvEVEcxaAmzrxfD/kxhuEHjPMFecRM7vQLAPcrnFYYmAHyi2GE8P5of8R4oo9v
wWu53fGwyCjldEJ4olsPjPdiS/zp9YY8VrRAnXDkcSs8Bd/Si4KpLv94ecl0UfRC
pIVAUOtlf/RSMidDOWYxi158ZuEV9uprHBSWWma6jhyRoAZIPke9wB7McHjCbm55
FeGOOYZqfUJs6fjnFW/22YsCx36yf2S6onmDxX/WEisqFp8nYWvaWL0GUoIc56ZT
EELQbHKe5/pIUNr3xlKN4ereRzCbeE/Go7MDm5ytQ/YFRMQ2O3Mkv08HTEXjmSft
66V3frgtuDpwXIAQWpNbUv9cCsXl1Ap708uZe0EqUFbOiDBtv3oPojZN18/i722h
Cf96bNqaescpLB04Z7Xc4BZDcNXql4eYCsv9+Lm8mglnC4+slx1oIoTPqIyVtzXs
TvxbCLGnElZH2MLCkaJPfW5tCcY6inOPVgAjbXVc+jX4UEf5EfE6YaT7faKqToTB
BUjyBrlwh7vX5ndyuW8cloe2AcvDClH1zz/G2LCkZvuBwD4AdW9UTWX8QGa/CbsI
HyLUrhydprCrXyOmZiXXDm7vIBZFwVX5RhVon6UDMLiNCRL0iXfOOJGbdpe+GrVA
KOOdCGY08jDVbzzjyTY/VTjlDv+AagRU7D/8whtwXqv/huulv3nKrhs6u0OduHzo
vJG5C6ecT6SeiyRUc+4yjdvOJuWk4UINnNwXy0UddE8t93ZcUlWY5Ejr+0j3AAqe
EuEg94+ftk+K6gS7GugSxlkrLg1pY7x+rVglD9i76+XgdzIMrNBaviA8UTWZoy6O
z6Y5B42rFLx0Cx28pntokR8uaFkDyeujArnrZQ+77Y34/3ufr+m0b3BNNwwIDP0w
R0YdpcyO4i9Sn0P3AYmVbcPUbtUNY4CMUsK3ymu+TexL+6JLMxvXDbGpgaaeA1sc
psVGk+ZY5j0eJXQJBSkyeRTW8Wa8tPsJaf0uTdFC0ZNTlTDkwJ2LMdItFGC4zpmt
PLSiZl3pJ/emM/+1se+RC+cyiaPogxS0euM77O3BXMpawVL2UO0+Ol9yJCJOlQKH
M+ga+tYNXVUQ+PXgl33sSEHG09yp4BQqJwrGsmeBa6/oWekJwxVYB6Hxm8cdgmBs
xf8s/SsvX5yIBhzlj4OzaTPfLDTO+LUHDNLmmcsQqVeoWst6pciePWx4IQKv2aKA
d3wNmd3ywfU1NFDHKm3XUcnLn/iCUz06eAVH3bjTxsomQVAhmkmZqKHxnXIXVcCV
pd6Gbt4A38IT+TK6QJFrvFUs2Xdi6HPhDBNBguV88jZpvgMeHfLMFESxtnOLxseD
4jq8ydbjw0zb5jOT/rVDgu2AQsuDl/8fD4jbzb+LcNl9b83zUz9ElISGRut/m8t7
7mniaEwVGBKXe9djVf5Tgix64Ljm2vOiejLvX4toj7jiqB0bDUPChOCRpZFPEEK1
W7iZ0696hJroMnWX2bZ+ILtN8X+i0cSmCQ0sd+c8M5BmraxquxGNHWk1D9l9nDBK
89h987nYDA09GvLvwxNDDeAG2BSy9dJBZ/D8B270mKh+Oqv7QHCTDXZQwJPI1Mvq
3A41P7+SUs9VvHFXxWCpDRINHmyV8GczfINTX2Y33ATs03k847WtPrfOiMOMS4kZ
NfcBnKrnWVRT3r+rXK3sE/OZ5jKMqWH4gRPlpF4tyijl2dQyuzD8zduxox8jhkGI
evNkcDTVbR0w41EKuFCiVeWffJNtJjzCnBlMAKpZCc6VjWIblNdUVNAb0LIadNrJ
c2pzRVy+H/iUxv92/kEZ4rwVBkjHRW5kRxyhXdUWaxImT3hWmVFBs1J/vTG1VbG8
eKj8yqTy2cWDCsLEp+h1u9a/VlfSqQuy/8KQTT/pXJML2mcAtIk94P+7jt49oSek
zS99IVG+iTxSK5AjVmxQSzauyXaZ+XjTjq0hjjhh2fsCpvlJngeSUmRSjLRdnTzl
qhxlXR85XUwZ0moj5V7dSfuoBEFhnsp+tnrOaAQAPksP6E88q5cpi0u1nWL9qqjw
rNb9ruWgMQgZMjJhyyGkFO4BX9jKy/LAnqOqWEPJbFCH4Qx05LIsmHSfgIh0ycwD
ZgQHw7ZxX1M33MvyOZ9V37NDW2OKP0xHWq1z5tq1JelyLRygd5BwZajUQie7hYn9
ZMLre7WUkX3OuHj+Z1a1UuVDXq0zHfjUrxNkI3mmN9Q8Y2gNmqDMuMa9g25CS2h7
A/Ug47n6TxhtFAXivCeyZWtX7Vp/B/Yf42kx/mRrI/pIj5ZNMU/9ZLrAtACJaMmt
D0pnifgpQlTgbouMTzU0YgB4WHOUi2wL1484pcd/8t06UtqL9CTScEllxTYQnyua
5Vc9kMi/scy/zbCDz9Vl0DqAvxXkSRZraQmuD3kulD23Z/fQwuoenEGgO4FrJkeP
rp2VAHvcg9edmeeU3tT5yK0THXWkcC1ppad6MUmZmQLGipEP0Tb2PErH7QnwdCjj
NjfBcRyNEDFXTyPdmX/2ImHL4kj28/4HBK0ZMBzuxT3c50/AtMqYxFP9UOixziIP
ZyerhmxLT25kJTr4o+IwhjNIg7KPiJ+Ji8Iu1vVIWq6W7jmjtSUerAvz3FnWGzh2
WX74p3UHfvxcuYB9aXVGSrhXCLwQMCZHYjcdIUvsFwuaXhQjV0pdXYoqvRJwQhiJ
68LLa0Ee+fgHGaKN8M7dpYFREBwK2w5ZDfpwKs113s+9r3c72iX2pn3gM1y8a559
KVN6iEcUx3uSXmaUJu+QDNBaBjxyD+SlRLEuXarUHZKxPqOOAHFj/Z/3WLE5a8wC
+F50XiNIYEMSeCDknG4PdEQ8R0EGrL9AIyBgj/YYabRhCABhpxXf0MSHkDQEWRUI
CB0BUESOuPXaRUF2ciToEvkiybSL4B54UijdHbM4HUxOvQ2NfPDY9/VWk1Qt3DtY
9sFKX2JtsH5lkpI2efqWzHUbqI9YXFVNGSyEts1CAvBpX6PtnZZ0f+1OenICZ4jp
XDNW5qr4FEGh9nZ04+Q46uu/D+yoRCRe17AzkRE2by5I6Lg07BXu3LVp5vUffoBJ
sUWJN4d1t91ezdJtXE7rgyMP+smfUqnBcU7/GMX+AY1G8sRd1SKjguKHqNeg8Duy
t1xnrGY/KYhbXPrKFm+a4pNqN9yAKaMy2ooFtNfkyOP4uWh3rqOJtio099CxeMHs
PkLiOKAAsJ/qb4yh5GeDfD5f/6fsj/8SPoy/cFOufQ9zUwRlfR3wIKagZcrui2ds
HEoEqoVk6f6fTeXICGHZfprzY1uJbA+Ql+9Mhz4cENP1TjSzrYgiiKBt1BrydHsT
p7samxQLtjJUTSPj6Ky4hXQe1cacGMtQ59G1C9RHh/ZotBDqG55+VseIdxk0ahAp
pNWgK4CmATEkoGH4dgc/F12Iau1GAUv6rRb/3aEKzrCMbU2muOrW4nh2rFs+ASlj
anCdb5h4sTHHmaQ2NaQiCDgKzNjncdGK0UGVQ/C+NFq3eB3sbeskTKU0VX5AH+mO
ARDjiLcshPq3Oe5TocwwJ64gKTdtl/VIgF55PqRwG7SwP7amn4umrtNMRk/ZXXha
ZloeMYIo6r7OwLksHc+cI4Lc6qWfUf7/pSLg++wK29DImxCzSogvU0haGCTnRflf
zHkMU6rNLwUXCKtZqGlN2GkjIzelwZ8rHPOpHn4BSTx+8kUo6w37wq3L5cB+Ap2g
DPSVasUC1lzd0Wd0ewMViEYasUxe6bUj0ojo9exylYE/rQTybHvnBLXBOXz7ECnD
lspvnMhl0mca2YeEuEGVELXxVOXtpUguDqMjfpbg3J9fn8Gm0dKtiW4BOROWHrBv
WZH/UbSgTNamHAjrJug/mANv4JNZLpsZx41JIc6PsQZAbztKpRRxvP6LH4ko/Kvj
xTE6qYJNLpb5Igot6D2A3FU9hJOFVcNf7TtxXdf5zgv8+Pt/7kOOuHR5AB8ZIkkY
/CsSToFE2Tot7Lbh6XaXL0ZWwN+YwynsKr8IuIDfb1invFm08wYWK4tA8IE52Sqs
T2flhWNIyy74VjAux/mbYiyMu0A37yGXy7/qsKUBaIrTlEB3xN4zdFqVMny7vCWc
c9fo3SGsPHaj6F3vMVTS+k0XnOB6bTcYxMD6teP5B/NfAtZbZ5TT6wVNZnZLIdl0
HyI8jNngwGMLvuaa72PaqWhYOcQzs4yxRQiEgd6s+h3WOyKFi4RYCJrNhL+oKAc/
4GCx57O9RMHsrVhu0CaHMd0GNEulOSd5aYF3EX/fumaK41pJbIz5SB44iaOA8TLF
NQoXEO6li0IBdl1ZC8PuV76GVcfkqNIxC3AfQ0uK7THa25y10Z/YXOLBhI+vA7d+
dn2A3fiLH/SsXmve2yh4X04C9ziEjgCUJ+xSbxn2s/rgjCV4HlNvDotG3K96hVLK
7KrdzmvpBbv2etQwZivyrvTqD/jwEWHtJgW8lJ7ywMOTa++GlzDV1I+coZ7iKwa5
YYMg0lWpZHeXeER2ZY4s+f9vfYk4pvYCYDeJH8oKsve/4wbESr6CJmxcz3T+tNqI
jQeBZj1ohzc9dRXeOEadMNj9vm+xvq6CyxY+3IKTeTuQ1XCVagoP0UCB6QjXlZk/
pdAmVmCjXojrYdvjQ4I0IgNnoXjbJ3OkMlzzUeHEVmUz0+Sz3/g+ydVSwQ34WZic
CjFZ4xByq+1p0t6AfRfzAhFVwrmLtdJmbKmfyPv7apMJZgb7IiFQGdcg6U1vIqaM
RzwsD8EVTENt3cyzVjSuWdxmSFqbNQ/j4xOSeJ2mrH7kAtcVjbdhpMCuBj7Lf53d
z8SUoOh2anH4goYkcAD9Mgbz84+8tMvZs6oG9sy6NDUPfezNZg4oUHjNMJduSY6c
8P9TOlHHQhe8XvfdZr7bauCb2mVU4LNDnHNPmX79S80IcNjacH3iHZ5+omEZVh6A
EexMz17V4w8oFq1wF3bhLtp0ZgQl2N/+8bLrDyP0kdv58/fJ2QS4gKCuCeOWwSCh
UJvOw6odwyBQ1csdaU4vpTHyqTEwcfWBdBYG6pC80HEfqmRVtYA6d9gkfwFI1bT3
/YGWRZXQU4JnzOrsUXRk7yBb+NUJMcUKHMYjxDVryvgQXPgoxdEZOlIHM3ycb2tS
X36pyZ4yoKsDOO7aElYJJxJjjxMRWNYirE2uFnp7J+21y4FnozzPUohFclHR9hyY
e38P5Vfu9pnPszLWOKIk81iPSMnLdBZShvEVL7s+aDJV6eTGhWstoN0s4E50xOb1
EycPSW+QD5UQdCbiyOS4PIQ5NxNfeCdzX9ixM7/ygTQyYYckK/GnwZxZMsolRlW4
+KC3SuSDvRdcYkOMd4QDFnmP1zBj9XWFc0HdZuiRjIZn3JGfDOshrw02+FCtDSMs
1dSeg8nLunehohsuE66E5WRfSqGrxP36ydm8ANAMd1zT67JVRWPCEnpYIupp178H
f4uXjnNAn73BoQjYKi5y8FAbkzE7w89hSQlvtQhkBmmku9tJtCON8XO7YO0k6gJ8
jmaVzvUWGFowCH0fyN4/qGxc5dmwIQCvGw40nutP85w/94Geh/0+fd0oLctGNtNU
xEHUPrc4B2bzVXXRchOXghNUBZo9kVtzwWN0iCjkfownYLPLabLG5rKOYkcvBFQz
QShrXEZq1X6iodnG6PxlT+4z4gzQNeqe6GarVKOlk0QVfEBB51O2fbGlBASLfJ0V
aC5JhEoiiYsO/bZklYWpszUOuzJq4K7Ft6khV9KEB1bsN31u853TWyQV7+2ViF+S
KfCt3q+tPhWjGdp6EmfTsPm8gksi22ZrM/K8mKj3r1g6AtbtCC6UWVLXnePjm/LA
tj/j3SmYQMTTegyCh5t/AVojf7CYrxlDmGVlRV34YeXdBoDL9HK2sx1CSYL9/Pug
FxmYOfmdtbB0G+ccZZaSmQcGRhVXjPZhC6bRoAPL6LA2Yv5gZaVPB5Dd+LLihTnm
Z3tSpjOJs4ONQsbshIjBKOGwZrXUuA5Nu1HTmcTPEB3yAR5HlO/oQIeyxZ6yhUHN
jSJnveD00TAnphN2jH88hrHwcLsVzxVhuwI+p1V+NoA+LETv74MiPKzRLuIX3gJS
c7jTebOp3CPQpfKDZyXMXsP3jNBF4lAFcxu/MJK1aO+qC79uNJguSBUD09rG8cEA
qHb5mjAXFhilBMgtzMHQuVp0uCFfttjYXfxzTuIFxOXsxif4oQf5M4ySamv3yFuI
EYvdD/5sPNcFEF4q9LbS7FTLNZnxr1Ulya4y8KnVEskrRoE6AC7VhffhULGViF0N
dP4zUhm/XJtX6tyDP1O29qbpA8IlQhr3dyj9eVDJQL4LPSzebi2wHQa48Q0t6m3s
TqvvYcT7OLYLAMEwp9qFZgSXDbdvQ0xa1PRf4vdOhudvb1r4MWev+ydLIfrp3Ru2
AQDc649kOw4w2/n+HOHxVskQhnZXytIdgN0MyUGh4sfXc7Ndg4AfPS36fUhW4Gvf
fNJgMERCJoezN0XrpBR+gn/wiUFWvCgtFaftcg8suAbeEGQgBZlHczAe69mG17BL
lpmEQhz4czGu8dMuglin0/DFRXLMsdMBmWqpIn5Ui4BbVZ1OwdbvP4ytB743kioZ
Z35IHodUsUkKhqgDQNNi/eqy18SW6dWeGKYKrpifJ5dfu3DcyImchnKNQecr1O2g
zy6C7sieOMVMNuEHOqefbniTQT2SyCkYvqKhj1J/KdT5RrA0eRz3ZbjEaMmk4fUQ
JJ1l3y5AiHsSRx3/XiS5k2aupT5KwIISSlz8KQ0/Vl/+Oh+rtwFcGr31C2RyufLL
8mf4YUUr5se6lAodkvpr2B+9/d/lifvNr6+k5XaaG3/forShnIBf0bMSFOvQmAEN
KQTVeVlgqFk/ZUWmU4zZA5HJzwlQpd7rbTuTr16R2elL6j7TpWwz3SuSwying8+Q
/JIXL0RT136YloOioSJ0QAeIRPVfIJgT2WCaTbZY1vq4ZKI0ncLtyNs6jTorRcC3
Rm5FqLEfBLk9byX2yyapxBUYrQuMlIXNM9/JSLwevFxBY6I5jPC1OkVTCc+nQptM
uX/bgSbE72wR3rlg5g29IpDLblhq+tRxVaJtTlCeIQhoIoGBEgFLaBYigZRDTKvg
NSBjJDumviCgTXnyom/ltXo/r06DLbHgosqhmgcGVavx5PDwW+Ix6LIjbfVv7DPL
Gb2TRmBl3uF9/9ZKxtX7S37ybMM+ZGyAUlMIVYb966yc6b1vhWTiVL4vXkTqZ2VW
Vq/97NM7FHWnH/ClKFr2Zes4xf/Cu0PCOgrbfbAf3DV+CxpgAZWoigDxdleIU08A
GmjJTuACrWwahWOvqSb3GSMnq9JFiOEZiT72X3wHsZTC/I/2/bzOOfu+a/TT4Xgp
MkGZAbdbj8BgGk2CqWXcIRClQRO1OxS9HA+GpPRlgYu1M9LKP2zlqH00qRZYMmFX
dV81Xe2Uun6L0h3VUIDgNBS00Uni/V+wkl7nddeHD3nDefJpbLdYtbHfEjrWbzuY
I1eQqNynlUL39ykKMNqnqe8l6/2PMLa4PJ+ERKjKDnBGMGeNxImN0AcI0qu+gIMP
xWNje/uDCzWg+cJ1DxwdGQDgZXx2kJgYI75yBD5bctvaXFmmL0MLtpvoYduEKWMQ
2AL7huk4dBTpsB6sl051nAFAYO+OTdOX45OSyGSG+Cvkzp3/N9Tr2lHO4vfwmPFn
HA6rmGP95BfhanlPtY0dqCTAF/61MZD5Im0zOdkDlWEP9lWOOeg/KTsXXdM6n01E
aqgKuJ7Z+DDpxTVb+2e70KJ4XLZ+2KGLjAFOM6VDsSnSGPw+wQAKTQaSDZDZCHIk
yiSjHdez/ixJ7xpUNp73Bmtf4TbJgP+ff20k2h6jpFvG95FqLtPVcEg51NS4OdzY
z5bP7A+TunHZ016hbJQpfeuokSxIKmTrj9giA5DRrwuEX6UKP5KP5nl8EXYeew/R
DH6ZvaSiDNVV4O2p9w5Zfj+YZyBuVvRsoFdsux5AjJuHYqhzh8CCFL4Np5Jr+90S
x2lI7fHI01AYamvQ378gmqi8usNoZGKIj3SLKpzNx23+Kpee4Kx5JUFKfoBeHrud
tPW9P1eFOGMG4JDRgIJOseLmeqwy8JhJg4XPXB4VbFyBQtLZbiml+K+4F1CC2JIa
+inP3n3dS4Ge0gHWQR8x4ccgRu7BwavGMLywoSqdO/kNzreAA9Fyo+Vei4MxjFNZ
c/0n2JntTAXE2HkYI1+ZG/f6l2MPBk8FDH39wifaISbvfNcS1VBf2HU4PZRr3e/A
9KgJX3hHOjjPySt2GwmVlGDg0E6KeNKYnScF4lZwg/PPsoyCQbZsnjF4co6HZkAv
1xurufykWReRZkUJg8n0HYPkVN5IwUFYyqgBHyPtnhyfHkH++6K75XdaAKX/z6ms
zyZDwT8mLWyRoyNPFUvc0YgbWL/yzshNJ76+wjIbKchXyg8TD6XXa0nG6I6EjSHk
JdlA4JnGR3Qlde11XBYNmxtrTnVekiEPKg55mPbTg6lrHW5f1zqnfDpvGzAuVjfL
EJkWKMZktuRqoyvHJZPaAPpZPdljwjlXhiqK/yr6XANu3pQiemaHWDNY0X1uaXN0
zUC//1YBCanp0PieVTWMZEN+6pmFIBTbRjCpJ7m6K47va21zwnrdLVmKIacm/kqD
XGHmsR+mlhstoiX5kEkNQJIX3Oi0W3xSWzm4Sl5Q46RFuz4ti7oYRchK7mEw+T8l
IMCvbjGNkOalCwUBOM3uECK6HaTEipQjdvsN/Zcu91KY+e4D9aOSATUJ+O2kebxV
FPybsiR5QEK6ntKEWHMUT1ix+vO02OCibh2z+zFN5cWMc5BPqinSvlKONuHecgZs
jVTWxvptVR/UIneeUO9VQUkbaL5nouUqQrXNGNT3y0uhh4/Nb6tUH+nU1wvTpJOk
1C5bbKjmUQ0ioXhVo9n6lxbglUBfGWByhc+kBijqXfIesBosfmYIW0e8LtZDUW4f
Jo16SH21QlMv+/DR9vzH5TpZ0nlm48BZ7XawglKfnZFO6PbfnkGokIuSIAwJwXib
pwbr/bLb+eeSn5Mfi3j6lUyGhUJ70/3MLeD4Ov4rDzdSrKveGbSEvSoENhKpOPAP
ynWBI2lXUXTQtQsG4BIjyo8IhmbASufB261zJNzN0qnlfC5KwPM3gAcwrPEOKHSe
EQw5nwQfRTKWF/5/NtZxa4D4myO2pTPaH4wpc0b2WdECFNs/ePw6VXaXxWzsa1an
DFpQFOOnqPVONJzzPqL8MBWfASKB2U3yR/XMbYr4nkqEkbNPfVHDINo5Qn/NaSQg
yjc0Mws4XWLQY4ZWW2HsGRo3JWiU0Y+Kl/UwbS682BgNkvoGlEEcfSIsedN9pEtB
K3XB7VIaSSphLcBJdEEzw7gcjQbgzpkHkhfDJRJm8sLfywH4t9RIB8fBlGAIjmaZ
KXbG5Fa5Tw+espmeJum8GgIT918NhkSvBMfTOY4q3qlXKJC1VsLEFH9zeqE1cdmZ
Sbo3YZmlNYlUntRlzaiYdnkZrQbZsF28iR+NdS85zXuNdxhnv0YTY6ysuQEemBOs
wna5dG51C55QjVplSk6DAn4ibtJh6ePtA8MU2+EyaRBrkx4TlQubCQ6DXwcnI43c
zm9zNOswGQSSk8paHx5Q+KUc5/NFbOA5i2Ie0D7hDAkVu3fWlOLXjEFgDUF48nWY
FgG8kcRuUycaSgz4/8J6Dc5f+CbotCn72GJsCyCvzkDSJr+IcDhgPObcgbXXBs9S
c14w0TrcGa40OXOY5BbxxiDFuw5TNgcEWOKqlVrkSWB3fjM223J7yylTu56G4EhX
bcBqqpCszwSYySKA/lZ/U24N0IF7djSkaGKaANHTk1Vy7aGg0lXDQToXgPUF91NW
yF4NddU1R759nhC7MIWUIEQISh9/H6Gfdz9OeXynhwRoOaeDdypVCHqo0LaC4MnR
lEsbv24d/Z/deCmp6Q8dIFLSkUU9yMv++E/tqOkQLbvOp5XK9ERyF5zvdn4wz4Ki
OqWxcJXX2LL3DqgEYnAQVSdaWfX9f4C/zkoF6IvT0ftLE5eCTDyRXwkJiRIYj4FH
El3YMFPmZxmed+OgZtHs6YTkCsVwblKe13/XiNAnheemsqAJ4kK+hN6CMfJRxkWb
On7Dn5BX581t8RUAYGBllKcr18S1FMAxAaPIQ3+81pZeC20RJwaAUW5KfKdsS1Rk
euW2WqUa7mRiuqmuzuZNiShk1GqGRJB1uHdT5cUsVWfs5p9G1ImKwIPcGvY7ykIg
blaAb4m7Ki4+wx6EDYyi4Gptwjypcq981Y0FTTFyH1XAKi0x0o+o9CrlQM1l7xjS
+1CrQPXU/Bl/SXebFkXhwzNNC/DGshTJ3MLFrAKhOCgVj4oEp0l115AKxpjR1msQ
V2Q946QVqYi632TPy1kY8wvUI8sDqgyet2RXhDc4d/rFxtKNsLfV8TLLvPiwYBzi
bR/dyL6RNeB4cZpsyQq7VZtPfQ380i0EyoO8mrWRHkT7raBAJJHS9naxh8B5tlQ5
Mb5KqzigMnPz+SeAehNXfqXE5VynnF1mgsrz/Y5Psr5ufhS0lEjWUm+LAd+jBtoG
C45sVeQV1ERu9aJ/2VGOa0tz3u0gFGK4vW+NCNrxjhyq0FI3diDtv8AvkjnZIa6I
gtbfJsNgpgW7qwedjoANNr+5lV5Sk2ZdR8mvlQo/w8TDhUFmWzIG4rNrcrs2+3ub
di0FJmxjEBqiKWGERap50zidNcsO/rO5xurrLTjjPG4CNy5CFvAE1vq4Zhca1WA7
txMeUFrcgg7otTFx7bGoNGoo+owzLUdmVZGLeRpOxQRLHc44QjU6ZeGcsfCq8zdC
q48IB6hH8OL/ETJuO6dZPUmMVohNbeC96ndlMd37IVnI0xADTQZ/zlhgbjOdH1tb
wLtQC1sK5ZJWnjJw3eLgG1EgjJOCLX3sMrfel5+5cXVdnAbrh3kCW1cfluJQfL9K
gNLGrZCvjaywyGVgtWja8HdMTZOFLE5TGe+mNxfFhIcP2vkPZ2llyUCkWBPFIkZe
/lILisXQAt6iPxLiDhx4tmjQlPk+Z6hqT2uz59w+rjIM1S4cw/kqbJdX8YxI4+Wj
a4rQeYCAUTLhAQxYxNwrDQ4UkA488xGkWeDg7uO8porTVjNQC6+iOzIdkfLggcO8
++hvDjsGyuLHFa/BvAeJOcktg/SHtqx8yM9DtIjUIEpfJf1j1uDMAFrs6pm3QLKU
HhQR91FwFRIug1KGoJAorKGjG9ohryDkWwCvV7ogWX3ub+ckMD4BT9jqIKPh6VI6
wRDxqD3sAu8bW6TUQvnV15UkNueaTLXHWFsFQ+VRUkgutkByylf97lI7O/T/9soy
bLsF8rUq8K50gauQRB6RbHNhelbaU6ht1k0P+DIhDUimR9oDOgpoDnzZzQc168SF
FT8J2NQTh/Xjv7mDUS3eI6cPkObw5FtB/2cgI7Yc62KUXUVhq637Kc4S0dfdW/+A
Z0ORLRFPo+aHeL3ii9PhORksnpk4lLmsMJ0uco056k60/tzdAk8k3Dy4CeHp4eOx
uzvYc1rehfi/jIs3ax282eY3+s4RpvaF9g9v93oQJNCD5FqG7kja2TqH4She+Drn
QSVY3HGWhvHRm9TiWNLOc9XZG5nFabJ8nctps/0yQWOvV0lqSEkVrXt+0+74KlbY
RUg4SVIfqNj/Sb6Smmlb1+cGXbzwwIeuXfCvn6t9fhdmSOw1enAXJ3zn2dXl35Fx
2C70BDZ7TTU8qZ+D9uVVnGjAMlJHYc2RhuRPVl8nnoVij/QIrPfLxkC23ZjExzmt
umXbh0Dww+ytq4VsDb6e+Wl2qXlOgFLKU5RV2MHtzTBuhbrF49d1NBtiucNjeJ0K
rNplIUcxUpIyNVbp3TWkeMyzr+ypaT6aA1nXqAvnRnhsmKhcU+yhk7EnOfSu52h8
9rfg5wAAdxcMG/Y5olxnDBUe9K4zk//P+vpXBeVMo7sBqxY28+jywZOdHoiUuM8t
XZhKVAH2V789j3ge9VLtgKy0gElcIwNTf90wtJUIpY4DE1kx+jODelQaMABvT+7A
X5UePUsB4qpOO8HHdjr1fKGfhEUb0vZmxm23B6vNE9PZqeyvlUqbzY2TIRc9joJj
x1UFHWcg8oy/ekkJ9E4/bpUBktBOJJzshx0JAUCFMebKLcb2lkCcsoGDt1ryTIMU
W9LENCNIlCu0PGWy1xblnEOh2VoJPITz4xej3zjBGD9EKUCfxM7UXjiF+GpDI5FK
qxeN5HgTrFNfRyA9vRlDHCKndoGvSlSbwxqlL2LjQZ2ininscQzVUTMQVz2YiG8w
j+83Hmb8egm5Hu+vvaDIkC+tmBn3L16AKqSKzYQ+ZtWJIXKkvio+iNXhjycQTibC
dki/m+sxlp3ICRM3afvuq84rAc4mPS07IWUWNBV8Om/1V1xROlIaEQc/ueQ0HhFC
VsBjxdhZcaZ6BKzeIRS5/ynLo+LvZrM3FcDpfwd9QZ1xLXeoXUwF4wWayFpjwDUm
4SZiKp5qEADR2rKSwk/B+Wg7BdKVQdipbojPVnFnXtEVgv4/MQ8441w2Nv4lVSts
O93gmUMwjTtA5l01B9Gp5BQ5+GCN7eiUiKdpRLQ3O4TZXqM+Z5+PY6vpP2ADvnoL
QWhtxZUo2JhpzPi+YjBgxFjPbZk4VH4nI4JbpOsK06JIMzQcjgBwJ+DTMOxQwaCs
rBaUK4anMG2CbvK0N3nF4x84wWpkBQz6Su1CW2d2OOQuVfIR92s6ExzfoOLh2772
9PyhVfo7n7UnKCHyezPHSzcXKhDn2DoSVFeAEi1sn/ud7167ibs0DhhxjiRRrvmO
uG7iqqO4I9jcB+pcXWtAsEdrZIlE6UcG3MWajH3ZAdFw/sllQ7jLYjKRIv4VmKz6
kwcqst+u/1gTH8HSJlB7LQ+7ACzFVJTI6ARLU7xX63zaphHsMh+4iwjNvFntDyKD
Hi0RGPYRWvSII2eg4pPxPdxlNt51eTm0ccJGjipSIasxeAXm+upjvfy0kaBrehlz
rFv7Z3xOsz9C1Gi2sBvt9SdWTEKPKMqDVCXggcoFpnZc7+BSQor1lGfdpY+hqR7V
ZoZz+0wq816nqO7VxI6MVjiQkZx4vEyXEoBgP32Iu3j1i/po+ScEhNrlswdvsHrO
2f7PXVlEZF2LYk0mwRnEZxYypu3f/iwKBJ2WKn8M401WaWk2kWoBpBxR/tbz6KqV
ORr9hbKDp+tJ69n/frPICiixa+/C4x+AW7bV48WXXqZclh6y+/rqvPzGe6iLzSGZ
unlitUDeIEiHsFKkYzZS0Eaj1ruMjbb716dXBS+G5apTnXIA5FX06+PdrcbDdzJk
np4HTH6zwFwinFHVfbPxdrHyC3WZoTWa/24BiVnphvCbzgWH1245T7O44opAzeWL
iBaqmU2+KqHGzUO2a4+f/f84KJe81gPCAymrqADAX4MCtLpzFRgwjcxFFZQ2e8LX
mdZCoDTF7eO7/nXZ0OwSipL97aPARucN7tnHOWFM5zRFtjFMGuMHgXdfrWydJzVY
gQ3DuNT/3BKEU+XWuw24ojDCSYNcfjKon1JHQ+voqkE/VK9FpLNvaJB0k8G6HCES
bNAbmTfNkJJPXEJ6QYqhVhZNaaiORt9S5xXW4dfZImDJ7I50P2/iocXXzd9eJdGN
4jhDnsYJ4UXGswiFfoRnnVJIUtD9BQOcoXfAk82XCu+SxruVrDosQE66ksMZLuEC
7Cf2R+GWGYVfK/iL5mYS8HoEpKQW13HPkRAfAkTqbW3MPge6WTlbf4kUvm3j5ISg
/igvbHlMJTUW+mAOv9lNnY3eGtlgHuUc7bD69owsFniLnXYK679811/WLxR5iRrm
Yfef+8dA5Ys1WVtAQy7OIWpgp3Jwv4pj0g0L2CA/1xC4fR7B+QQJeLaO5dxVvowe
WcSciG4fbcGm2h8N06zipljCrGfOp0snlIqmQWDFfvdCjnNVZoU1nGvKtxCtefCP
6dSpsxPpWKS3uKHVGb5d4lQlVHhnMccm0QLMyozcRc9U4h2cip9xJOcVw+DVTzJd
3mO7UDNEnnVrXighAcJFWEB7UE4Ro5dmq76lQq3aL6KahtzReeiyYd/u2za1PRqE
pGcKYObniOoncE06V9kcQiPktoW+Iko72w3FMK2/+CrUbn0pAjWxH3ds7ahbOKZo
abjdfbTf2vZjU2aqRptoV2uTdpoc2FQi6Wt7KwQb3xYl7trkEXWbwEqs8geUo3XU
2PV9osl7qkP0gT0v0z4oWfaNMKNXxKm1n4Ms/dm1hOhT7xPyZ1w2RPJE9M88XTLN
ssuTiiqPwXIsDua5gwuK4YbD6YWd/hKRISCdYhqMxcko6hXY+5Bkxxo5/UA+t3eD
g/FHsd8PrrjYyvmTTI1IWUe3IfhUrvMzIn+98m98ayByfnx5X0nkEHba7NBOhOIO
LJWKGrC5vcRs6/OYdTIoEGFduVTN90O73Qqi8KQ4E7gNdFOXWtp3NwoBTM9S2fPb
x5N9Sunbb0a9OF5zatVnnfS/36Z03WWXMpLBs0tOnxPD3eKN5aZboVYakEJMXcKy
72dvWsZY/CMQAp5wlvF+cRTlRG3bmD+kAuUiRvh+02slsCkTnY2bINqlIVy1sUaA
PzsPW6I35PU0gA9x5zSemsyENM7fprGsJX0uzCauqg5O1a9M9dexWJdZ5L4UxcL/
oUT+Goui4sqedNpiPJO+L/Y+Z1tviwN957yJBJ2GXT2Ck/hhBkKNA5Le0XQL35kA
Gh48NTiB8UDkmUcPezyPi/XFKpHeoDLweK++TDOa6gQWQQVfsmCM4WcMsX9/V7WS
EZNwBKOxqfg5Gky0hU6hEulFoxVQF/s4LrECHTS3HA9qroWHnQEqnNHP0WOExL/a
cP+M43lqKYI0ENcqops8uD1oW60f6yt2VslE/8bUzEAtELM36nh03to+C4CRBD7g
o57pu6l8TRfrh0c+YNmMY0eyrZgn1y8AzJ15d0Y6tH7cB5pnk99fTnTxx362exy2
CxZaWKiOWDxdxX19U1YTdTn2h9S+SoEHykCiMO/xZYgSHK+LLTazCxbPyJQq2h3k
Hh5aKQObgpI5+yDKNWiCtmHjOUE1UKOPMeVqrLa7S5o4+egnDhtVYpbT9bsQjTZI
QuIYgaU1ThSXKD7QIXmgkV/6gzcGK7kDfjUbLwpoIlxT3YCcLv9aTZ3pcLxZ3p5x
uKssnXPkCwg4yjRRPSYy0w8/C2qW+y9yQ7t0k9Xga7p6msSEgeSnt2pRwrPYtSC8
n4I/GvYLvCegWem6Ej9Mb92u/pdnWXmuJZudNPjDxOM1zzntoJvRx7GHV58D+oYR
LXeazdTiQ1Loj+BIe5kbRbuqR/hoczO5GfkAxswCnpTfk9axNPZsiy/WgZS2NU3H
UG2qH2xcjMg2bxdBRHfEK1qQ07G6kvTQ9R/p/Nre1sfsm9W+uGmDvnL3zdOpOv55
dYbuaVsJTAhLmmEc6F4SzxTKRsPfmakuD5wA4ECnDqng1X8LZZAOwaSZ16gcpzmx
y43spTBq7yvUixH6bZGGb0W0aTR5llQgprA//7NQhk5geC8aYq+cwT1aZZ1D1/3V
DJon5L0B2972Oql7EwYY0pmBH7wVcBnxWSSCpX+LjL4vsOByN373wGYzyec9OuPl
IzW+K0wh/hw9PbhqBrAbcPHS2AJmcp2TnKcGVOdhmW44C5H5ML5mmVwICFAHNvOH
hnYVAFvMTDYPIW5bWRljb920S0h4YdNbPud4TNv4O2wWkvJvp5eZ4A9rc8woB/5m
8OYdCNx/0WlrRSqE7emZt7BqVfiSa+zuvhMZs/J7Mq6ddDLrO/m7CQvNYkmHcUzM
xJxvnX9NO2YG7ivhQBlnwkqB4HTxHv2/UzW1py4CD7XAAlZUTIu/8mF/toJU7/LS
gIaGpbA4sPopcSeJ4SP+Ja9eDhqmktBTHD/VzgnTr8Eyd0hHAaKuDf44Rzn5s2q2
sk9myiVV/K00yvlLlpYS3TAjzvg4RgeGC+0WJiwwI9bZ5NolqYt+WRk8yyEmrnEB
kCKYIxORTDdHpBEE4KMaOctcqYetbYGKrllwWVI660j0CyUH+kTvGklajF82TW30
XTfakcEXiw9d9+72kZ42kZ6uFCOBYJHPbdZoQtB3rurz+bYqRAWYuNK9qr8HAz7S
7JHlx004jmPMkp7vU8vUrb+uV5+FqOtDcVIRBc9mja8EIbuE4CCPF/srfmKhIEPN
I5UG6pwPIwHqEVWG+gdn6532UPG2Nw02zNFc4dIYMKIRM9zMYaxc+mT1CkBtUcjG
rPqbUXV46fWZYHsboyxfjqcBD5kgzzrvuOgnv+/UDwJQ7/LWzCD780na/sbmaZXh
/FAkyOI3tc/U+lPprqlSL/k3s0okYyktrXzoe1qa5Xm45qi0tnTaxOD6ZbTRwj9T
xT3e01yfa3ZY1JUMO9IDDZmWA/znJMofr+bMvakFBAkZGiVrIOH5srFe1WZpX9RX
XY9Pq8okeQRJK8YJlZjARkTmxK/DTF6fOvAjHhHUzzDZuZ9G+McZsAxgBDYM8FAP
egotftop25KqjLBIgI9I6B3BBjZeH9CRO6VfQUlIDtXPwxI4b0vVv+mWq76nm5c0
FxNzKl2P14xnsO4gDj5KX+nGLB3nbIE6T/KYYtee+dmIMo4ldrzbQTrFNwWDSusO
idb/eaE9GJKtFABblcAfzPo8AKAHxuyDJ/vpe3WfY98GdBCwJQxqbOy+KacYV58J
Jp74y7NT6CMsg7kP3VsFSPUwc+Zyn8JJvmnVv8pATSwC3CGju/NIQgrdxzyjIlV2
BZxe9cK+3kzsV2vYJF9f/FeKPwvUXaJey+iS1g1EfTL1ElzyvBIw6qRvgTd4Lt9/
2lA5CWsakJU5ZG/hjPDi1B/bZt1reA1flhE8agEZi6bpgwtX7pshAOb5CbxpwvmL
5yQoilE4Ip05s3aMW8XObNaggVqAYp4QmzLy9+ZSfUVPaq/AKK8qt0e9ZDLn7et6
3AMxrHFLKo3VqMzI2/5eGPkgFdMJAHPYEaaayS/Q9r/NkSffUt9kdFyrlmDjph4M
XWEBTRDGJu5soVUForqKIgwwtMox8eCpHFZVpolCbK8Ng0dbcFbLpsu5ghCFEnxH
mwQ5fEcPwFimQbDR0gjvvKOlC6ZWwm07wbE38DF5rroD/yMQJmsQfHpxRWffhkza
IaOf//YyF/eDxBQ9JlSn4+j0HO7QBW2ppjg0kmbN9sT+bT0Thz1l9PiZxe9Eg6KW
9yoxUwRKB6HJQlkiuvWsB+3xNeXLFkiaBJ1yIvjdCds2VcQhlxJDJn0F3hcV6hha
ljMsIRHvIhra8J/ARK5mEE3BUl4/DlBPDGgtNihGgO+gbAnGU/vx//udhxHczWog
tKIeK35RfqUenYL3xvuWPN1Ef2HJBBMRIeq7eSJm+SUURrffgcm7IrYvrh1VNRcZ
EuZxna4WJmqOndUrG09AQxdO4W1iB6menz6yRE4FXjCPAOgWhkrkgGs54xDBUaTJ
6XcSuRQlk02kRU5zP/AbL3vCefTp7sSUFXs9vxAJGdS54Ma7PPKC4xJTLX11czzi
7xNdS6bVVolkSkZWL0B76Y/AQXt07+kyJdERR9vEYlAGX8DCJRybn5n+0P8atQ5G
Z+4mVhbFjjz3c+YL050PTfn9hUnjA/VD6lI19UYIxvMZOKQYqTVxtCNOc3SSQ2/x
5GJMS7mbVNTvYAn9cT7eqU7XdrByHQihinni/aOhdXOo5omC5unmJmEyOyF8gwoM
RbqgA2lP68X2/jKDNj0bpktYfpgUrr7amuVtp/9Du5mFFF2jEzyU0AoRXFQbFExc
SsBDJ3HItzABCDp2XkY5/h09Jojb+u6lEjeWNYqQ9wVMNUV/nSy88kTFnIAJ9cCx
2YDN3X8FodnxPX3ZbY9Iioh0NVAh68F3/2WplwVfTywND92V34fXf1gxMdFoD4kA
o1LzPOF/KSWrcnh3GjUmDY9FpiTkhWBW4g8GGo5r5JXSBvcSkCh05LKuA49p438v
LYtroyNb20cBcBkGd10XLkimV7B37wPu2R9HcMYQeYokaXUOMkes18H87SxOwD9o
zFEFoXWgtrdaDPe3KHNMzj55Li8tII8O2+xyGNAhB2v6RIrj6YHzPOzaKM7pCJf6
bFsDomhs48JZMl7hfgXNc+GtbJ6Po80AgSJR977gosO/JxrcDsOE4NgRF5iu+idp
Ix3vy0VYlLaFLPb5aSxkYjaI8VPQzKy3Z+is3OYOj/hU4UwRieYMXFbtj+XIJ3ST
aZ7qxqBjC9lBQStQqxofGQF4pQyUql0aJLzcxNMIiSEVRm/OYJ9UBgH3hCHVm7GS
3WeHQypUgjYlCZNzJlIba4fsoKeb1UEfFZO0Yzaw1hvJH7CNKOf8jWEAvlUODZ7a
tq2q6QBkcvPaUvza8uhk4CUrX7EsX88XN5GFSriNSHbefK4HnGuyi9pZhFpxFfGV
mcL7F+xdCdlH6Hm/4jlTKmxmrzPkQAsfOCBh5/bhLUSFBeo8zqXhFZl5KV/FRv6F
uJAKL6PzcifjVOzJiq3KfxDktWBD39lhqAkCg9DeSdRu9e8xszBgx85XoU6fOqNP
O2vWgN/HT/xX7zQr3MZk9iw9vbvWI5LDQAvsRIcILJndt2ixa9NGjADOQ454V9ld
cK/4dEGkCsj0gWNz3BCxOhksos4gIrvfmNZBQYYNnHDvod20aBI777jBZNi2FBZD
N8OZtGmdSR6+z8UYZSitI8Ve01fMypD/U+/I0tGOVIjBs74VcRWSA0YX3ICPlQpV
6FGLQt9Zo+Sh9h+1t292Ft9jLIEfDqWpRAB0gONwaE1GSR/EQESZM36YSDtOMIBR
1qQLfSCXfMORPv6NJG5RcmPQx2wQQBnqKUXnt1KL8jCHoRBl2vTTDFziiCA8Gf3Z
pgDdhyIMgtq6s+J887nfyHV+z4lP/H4gPLOj7R/Y3Uequa7iLcPW7UX+/ribvO/u
TXrd8neBLW5h7GQpeBBzsoO36TQ4T5eXp7Qqn0VtNOwDedw5ruBxWVTLAE2Om+Dr
xOaWf8KwUtzl/4avmo0zWrbkNdVssQXiUzr3h1y47ENznHzxdF/y0ILW3dhbtyOd
/WJRZC3UVjIjr7DalHBZgL138Dq2tLZBRPjQHXB8s42uqTx8754QCtoi3npq5y9S
19lhJWyMrBjJ36R0YFgpG4pMqeahzPadtZmWOO4n+eyVR7Txy0bAfFXwgELRm+Ea
dR68Y4gJVLLHiAmQM7pznzfr9kC2NzoO10KyM8t4n1GzZC8Z/gxfYLF48/mwIMUD
cbQGsaxxy+9bi8kxjUZY7xntLeUiofRWkk2/DTxBWy8EgzeLV9/2OU7i2YJ2tH+S
aRKYnZPRRKlcm1vkD9JaHLmBUwhSKt1i6DHcJ1oOrXkD0Lx7Dhf5VqCq7wrr/9cI
kWZ2V6rtvGrm0KBkl6sRx5KsNA8mVgPcerMsDDNw3YuPNmMZ2inG8+KEIIbZ996c
jSr+UE3zD2QpF+vHcfVC8ksLKjnJ8y/aNpjjYZf6KSiH1OrhPbK2wzLURcPgdggw
FPIR01nYO7cpraDqu7Yw5Kw0UN620rQQrSD/bH2PpfVVIMjA69yklqw6qMLuu+Tb
oo+Jkg2cI/Zj9HMr0RYxZLPnx+Q8P5xDVN4svenJNRfxCJjgDdY6+SSSd+70eDYn
psnBryZqdDJqsU3TUHUv4Vsbp/sh3TFzFtJEFpW16Ay0vIM2uPE7vdX3ACO3wCBF
6QUiIx8f9ieF8G10+pFw6JfQUvWrotG7Oi6X+fX9mXZMGpjzu50/M4QULd/oKvt3
Qxp7+0lbSA5OxTWWfCz9dFhCGszuJ1CGqHQ+0kQ8kUksVSqVecxC+/SNDvYny7I1
dxQc9vzRA2VY+tlpm1dKtJzXDnNvIJJs3a/A4nb4NfaoH+ww4eUh3Hy7JVusCDLt
wbd7Fqx40ntjyMV4fTwY55p5nOCMOCyJHw5OyTv4FP/qAJmKqZYTeVK2KVHTNPmO
Hv4+OjBqNaekLJq4pmudRZTyhwY0/uzTRuFY/ZD2X1ZNsmushcJcjcYr+1vUVCgz
IZBnOvz6BcTfSG5YT0JYL9vL8FDRHgc94v62ncqqQnb6SY9PxfQlTTk8GDyLkDPb
Q4dGjWi2sKFYpiEcF1oDZfOFXkwC/QCuoBFxYIlRzhLfeckLTztFa/QDhQRE9GpC
KOp6nb4tluIJZ/bUCDnxqEF/Laqf35UGVVtKhWjbJ6+7YvF7Z4QXn1tL24uja4pU
LChEIJd+WxuXwaUCsaH/QrVzE/oBHXASlUXiOk9vdzhXBs83p4bpedhttSifKiEO
iB0Jlci1f5s9xcwEQHCtYEhvqq5ynCWZL/dia3uCNBSUmedh64xLQw8pxjTSXhnM
xv5mO1MQHFnXqa7qQ57dLgSQAhQQTceqJTfWhgKf9hN8Rzvol7PsuqzkDNAJ5gtY
ParoaTJ3FTJTgEMqWpqw5Jnj/jd+ltHMXmoMuZiKhsYz1E7ojX2H38hz2sMnQjY7
L9WxJu/xUOmGM9xdIFQHypXKA/VtFyaVuX5eig3EkCo3ucqxDcTDiUt7dQfEGlnq
BGmofzljRD6KmzOgCQbWnT+tiHVLgW7bduXiglE8k6ZsuKFyZldsqpIHZVeSfphD
ItHk/H5rl1p8pG26syGNhsW9uvH1FW9dCGWYCrW1hZ8DPyzDcBnBUhFa99DOpBXl
qN12Sqqq1ffMzSaezWOAMi4xDJB9lxgEEn4q65ZZqV1S6T9G2FYGFmD3eKG2gZ9d
hTHLIHIqP7vze1UjsO2Rr0Y882rSnS/OBIjhHVE1KOzzk4DhvzeGbvyoE3RnCkRi
h4WqROAULXOfVZi5qWtcmqsDynQkiNwYeMkpAbqvqU4lSFtm1QWvrALStTnRCWJO
KMJb1QNlj/LFNOISlGbHBmwsjt8xhKTdruGucpDgJzykATBUR5TVGip11LvAOXpK
nmLT/wDooDKZlrl0mdkz3Gr06zBmn2h/geSY5NhbFiu1L24kQOJhBPi4MjOSk/ik
JNhKOajQwAxgyiEaE0MfA1ANBoUrCKSJkWsPp3rBhn+ySX+hdr0MJmpqQDS+18dr
9vCNf/MPpWipJSchDkYK8EKeGU5e9al8kRxQqLMke59CZcObw63HYi8QnVsmz37P
xxlvE5tnVfkUsCPj0UPTCzI2dzUgK62QV3NF/8TZCzZzeZLlJTa0OJ34x1xWmUjX
E1CdfK6PVzVhjdBaf2ZFU1DOzJZ6XrfwTBtSYUNsB7yhfxbOdYzitmTAbinx7ZiC
T6Vi+qA3Dd0xQzUBEIceVB8rFTIiOB7scSZWU4wpteUth0N3JtmW3V1wO3YaM6jo
Uw2/XMT3Rfo95j7xP+WPxYuG+m4H/LX3ELFBue+Z2944HYMQGrRl2Nzhz4211jrL
GPIKmbNCZe4j5bJz/CD/bK3qX+cPDpGaj/MrdDhPgqWoAo3pn8Vmap5btj/+o/v2
iFjE/jpEigl3fY7b0y+T6BXw16u/Ry2xAWgHURTyi+LEG9JvlQzBr5KlcjiLpFSd
GdcizMrPQ99yh5bj5jt3tgcNkKuPRtwIDMwfICXnHdKiUzW0s4kax0bqivm6pLiO
hHIfmaALB2Z1V3DZrgYJQN13UPGa7ABQqCJSnilW8FH2pRklHHGRXBLe3MPJmnJ7
T5uQACPfcomigw3VLYG0tyLlGr6QwX3GQ4YMcPEy9MPocsw69vhpWusMN+91utjS
lx/OiiHNaV3BZB0JvHDkL9lajGvlfJO2Y1FUsEEYPbJay++xoUD4dGX+V/0v0Y/3
72+oaidmgUeRMOQoPXbnK2oKv3E3VYq2oN6VphY8Gl90h2g0TEdYIFPPiAphu0J5
R62j6sTg/H8j3DYB1Ov7cT8yNzaeXQZjfhlXHxLCC8BEwrhcdkiuDZ/sqX76T5oq
hNARLv+gegTmQAP2/tM4E0/twVIynl4JyMJnpR9aix115DsDL0VyVz9ggO+uaogQ
2KaeX0Y4/FW9WxNricV27erxidIFs4FxXKHJwnsFNR30DslgKa3t3GbW9cMek7bH
8gdf1QQDnO1CQvbFVlwbyB9iAeg+3Ro2OdIvDjX63/jDR9QEICrM3IFbxjICNIKr
/bNRrlcvQ0RvGX60L/wunVrUK6P80SSIv2gNLWkXp3SI08Fm5SS/eIZdDH878j9A
cDhGgJ7/OYxeKjP48NCqLfx+Hgwd66a9sSDVY6/KHdUxm05Uv+h+LuJZYysWz22W
XVQu6TJQc1hxRZj4L5kfVUp5qTF0RBEAmMOwqE3Rp1wXWhIEHHCrCMnlH+wP6iZ6
nr/H3vp/OkLr4pCHa251a12guLIn3WlO4Fcnnpn59mIMt2aIAnh9iJUsXZ21N3bK
25dIYYOMUc+rF6J9W8r3Dg8Ocd8FRZZy0REE0HL8RRLQnmA+D0Bb2EjG/speoEXn
Y0auvS1JQFf+RZGPgo+lWWRaNCyR9bR5L0vvsGnTpttVwZh+dUxcpJqHuvFegKUf
gXEuVkwbKekxOf6boQG2Qv56UgQXohOwobhnD2k2TUvKhEb6StcxoTaDHaVRn5S3
sXt6m39aFS6Rq21OE3vy2CeADB1KF7cQVouVGSV32yK2jKb4o+nDeQUYQEMfq/aH
2ZVjLdLnYKUX9MsBQRyaN/gnsYE6Ywp2/8m/drvE1CEd+89PvmntQ70RS8pl7cJx
s08FMVmRUd8GFFWU6q1AuWFTvA5fk2CLQOGr0SEhEuRL01UJrLxI6Q6QERiavQr1
f6nAAuDXCe1/7wWK+4SYD/gmEzgBmCtKR0v5cIdlKItLYnEHA9+2QhRAy7XE/JBD
BFgtf1H9dyL7VW9LqLMzpsoE6jVy8ZGv4N4Qvmr+5w3uGLgbM2Ckcmpyxcm0rMbC
InMKiJqGrxhI/c6D+RFBuXjDzA7YOziWc0ygUXZhVjnWk35rAHup30IegwGcnA5P
hFJuf8Q3VSuNmAksoXcP704krk8Fjr3QtWpXCA4fl8v9/iNg4IyQv1wAoh89n/OF
YD5iUYSsvGhBlobI1er1pX49ulpuecsH8Vdj+d2/dXfDYxqNEeGVcTnRnbE8VHtz
1iVL9Z/zYuDcn5dJwwQbQBv/L402wWlxArQNb0A/3jSzvmmjXOaaUlzQscaDnx2n
OmmnYwfVrJj+BbMlnPAybajd/BnTTJt4eqsgEUrR8ZvHdr8dFoNMmvovMee0u99T
08o4MlEyj5f/pjfJ9pZBUbzOvZHUVf5QDmdjk734jpIEjBtYqIh0+E5wy4cu43eA
EL3b/opOhGYxhfiLIYw4/7nUTnH8TiOgKf5+m8H2VurqhGVd7kQTcYAHD/egLmg1
D5ZWcIcFEIS8f4wcZ8BlmE+HBWiWScrCQHcxxwPB2Rkdr8TkkF/jTGIcjC0u7Ls1
6+xfurohyd0tQMM+umTwqp0XFT/eIcSgm62QUuXtHkcCFFsS3jCJXmlo8IYF3WjM
MVhCo+NFQJfrq+rrJC1658M/ZljE7bFLeGRadN+6wGy6JotC10E1EsF49qxLNMDg
V+lbML3FL6BTMiC1PL8tYoojVFPsYdSq1GoR0/8cERZjEPPaNvAeE+4vNtcPLPJ8
suvRR0WhYtltVJ9DUpGQFGx/F0cc6FcVDObXrB3DpUj0NLSqrmvW08agNDaLIqjm
fa+3O5nptHfzz76+nnXYihXirJ97e+eu6FkfCLVwUdhJdqLCjWTdYvJuOfrmYnFk
TPkKBnT5f672UbivE64xfkZCh73tXtlBpGubCSxAM0Ex9P9yfTP7cuopWCVZ8ehc
r9C9IhuTzgbm/iLBi1tRGrDJPfjOCIDHpSsnujPO8+nha53+8l9XZfr7+ztbFrok
CNMDDGctSrU8ieUPXxJ33w5zpqaL4SMe2i+MkWBe2Cy/wM8JCva2m7yodKORFH0r
SeHZi2FSR49+WxCg5+t+G4NkSUxtMp3DfloZFxbi8RXs9shs/QLhr7Ep9Ruq0AiP
I0Y3YZpUjS/Bv1IotmV/kDHUU1W3cq7Y8XXJ/BCE9u5iHc23nTjnMVeRe+GJcofr
GRi/STGKWFT7+dw/hxBlrWdRH9zQ+V3RTn4p1SHMrjLCsXv7wQlmxoYLoHjb+5VO
h8j93aIQhtfCn6pmRo2FXLHDIMdF09Zy6tyrtMnAmUSVA5S+xUWY61bbv/PGcLlE
hkRWlpkb0+moDJq59M9L13Bg4GXwP7gSZi2tCpRmaWZ6yBCO8Ep7616egHT2fMKy
a6siQ4Oj3w1iwjs6TdyIJKKiorzac1EkGxxIJfhrPhlHmB5VVYqCB1lbqcNGKSR7
C+E+qzXx9aHYGG7Mj6dzyqCKZWP89+R1EjLHFvnnwGMYoC2fRnE/j0SYPZQTvTLu
68BP1ZwiCTNzObCRNmpFhVBNlrEOwXX52rtKh72KEPuUdUdbZLfzHSp3SbBdgL4U
vsbDbO4k1sYPFwrGHAmUVKIb2tFJ4u20O5+CTDAzfJOJ2c64Pn5WJHiuAjoY/6Oy
tuZDR8pU6T7Vh1tGtonFnHkwmyAPkaslTpetdcGDVfXFUfd7aoaUQew1tVmfIB7w
5saZdBEo1LjYGb97iNEZ9DuUPKnFAFl3oFnteoOmwbDBFfhTiyZ+dyz6pH1iURwJ
z/Cgmb10OOLl0B22WUKum6GlmV4ZE2iDCj6kPWiOgcctXbrBrbGsH+FJvKDEB74T
R3zVQ33dvX4pxp4cVU58GeINuOfgWXVyP2NqRK3v23HEZdxcli+iz3QfGl9/OB8D
U7+RXASGBBgUmfQI9wZiful6+8AlCOS3TPL+UjBx7tGU50REDT1nWOK/h5enT/v5
Jdl1SOnhW11Rwf60Xn13kIfKLEHnzcJx1SUY95CQlnaB1ZAiYTOFWmbdjA7Emj4q
WHA/SwEQ61VLkVwtbEHgZAaQAD4BgBk15JHCvf5d3xgcMiqkn+Eg5H/Z3UmtOM8n
29G/yluNmLTMALSNBLW9+fzvTJRQWewbN755/gAfLkexNISYZ+1tw7MYXKR3k901
uTCtebraacbC7YBDRuoHrQe7mb717VNiC+/3hYhdIb+pwebcjNYmsbGOqHCS+WHu
yAkuC1NmJuQT0rrmPO5eWo1vk+wv3nBkDcGA7CqvxouOwExEtOUTAoQKRS8oM6bv
EPTswGwGpdPZVnhXfEsYBkfWX+cQ3PLqbRnq/yuUei4rcPoQLxn9aDRSyHbpI6nw
L0Ky3i+4UIyTRCsid36qpZZxm6EugQmHLijhxZMNhQzUv6okziqO8SWLbyoC6o9G
OZOODcKr5yYDSgGGmOGA5kylKN8Q3vQLYvFt1nVpeez5+SjHFaNmahegQ5EHqWqy
vTa8Cayr30wI9Tap02hZoZ6mqYvZDtkg6nRF+7h/UkDWsKD+xMTsYVUhmuRmhAVC
Q0dPxFySV8WZP3y4rm3+2n8vNmXoPFRmqisPtUfHdMF4fyhTK8Tu0CbpspCOLj7L
C9z9dfThoxrfYUqoZfj2Z8n9PU0s/dLv04oahTs6cBqIbNXidnDHzAIysgyG2PgC
hBxT8RnyzZuXp7F+8J4BjCPLt6bks6yEH0PvI/h5rozNkud0Q4xCvgsSv8JWUOTG
hXkl8qdhIbBUi6i7En2i1MLV+gYrDIEaa6i5UB3+KlaP3VESHvlFWjG6y9xTUNLp
2VW8wOVfLh4xtXgjxU+0qXsMXtROXgx+PYqJgftTylVs/iFpKnzqG6gXSZNrBJwl
6aCcVXUZ0l+RTSAotpYscx+DjcedU0gv6PDddHCC2W/QYgm6YtSuUwBXuuPQTTd6
9XpkipkBJXuNuXeNknRheE0eLqQvnFPMymSTNjzIx/MsbPvamssoOG2+q3NkvDt7
n8umqyBrMNiWGwr1ORLakqSTdadLpYAfcN2MociHzMbmvrPVWZ8M38qmUqUQ3lDD
ziw6O9O4dBDdAUmiSuyi35QjUfjEJeUKQlpP30x+jI/k1lgx6qzq69Cue1Vic9oZ
dsJv8Wa33U5xrivpf+kKVNG/T0+j3hbPjvLHwwxxYi/y8xTsJeqzy9NAIQfrcAMf
6zGmmbqjK9BVMYDTFERJqbqzGJCPiiNzGTDWTmSZcaKuvtT/6p+qK3JOYolomjLn
keAZwuWOCGXryNSMR7eBovQjn4L88fnpBFjD4AWTmjXc12iWTtko6a6+fr+RGLvS
35zkqNH2lJpeCB1MKlLXaHYN3xn/Hu7YP62NIhrChM9YW57Owip7wsxaJ/WgJLjG
GoYObNlSYvyngCcoew9nP08okjFdt/T4tO7Cd7Ayb1OpRCRPZxfi/w4H0xLEXxVl
iUF7t9onfS07B0NM7SxbM1BwdUg01j22KAOFxl3cmIMHpvwTpWa6v39UAb4zwC8E
EYge+KnnzysgWTzPemb18ZJoyPwomXayRJ7WnouRAfjPvi5l/98f3farnoecrmh7
UXPQg/4H5nJvUpgjOpt/QoNT8rMKJ02uatuNgaRzjM9F4iPNTmrDkDC1dChg9UgX
0sc1wktWu9LYBU2fhNKTsMGjWwgI0o54trY3cb1MBx0WL9nKANoBBeFjjpBsYRPX
P98F91KAZ1TBaSieaF1TRpVz7zP04MGOaTJCvOHhHfmEPSop5Yz5DhGkLzYujA5H
fByx8XC2hWMZV+MHTkxPyrEhzST91qlr3xbuv+GsNMgeXERZTSeQHqX8LAzYnF5R
+WcDg6KjJz5MUQJT/5zR4ivjJMtyQIbNk1DhX3YdMQ5fvzFizBNYHlAsxl2v0C/g
Mnb/QSPOnoHYfttX1wfYtcPFNHiK2TCgAs6n1MSmo5kO4WmJ02PpS9FP2u4PIW7k
UwHB6LHqdxkzzXj9GZvhRz7cLOy/SEAGk1dfmNIydUg7lw+17SLPmohVSX3s8kuC
BL0NrFO0iFwMW7WBHBRv8Y1JpNSPag49R1omc4zCWmGmO+7/cC95l/80/XLLYs0n
DpW7FqLl+fNFVXZa7r+cgOnGUgfHTTnf+NXFf9ipp4ozNMwqJZvYtHWf5/ehj5cO
Y/HdIfyBnj/Zm8DbYJHYBFcSxnFbD3AnGfKDJcSTKKMVvAXpZc+lRkZ2tO42vczm
y6cy9+ouYxp+BQNUqadJsmhEKr3ZhvhOnglHVMrxr3TVxlUykfg7hpE4f1iir8t2
jQ+J40mVMCf8BEBPTdsAGG1Ngsf0zwXy66XK60/l03nDTIgSThIx4NRDDhwZf+Q8
vc1Be9OMPINySWpjcbTS0Oy80OdTeJYt7ge72wAoa4HevnH3xNNYfL6CXIq2N3La
Na+yx1qnhRZK4VpdXLgam0sC1eGkvCz0/fqXzDm1ck4A5lIGoeZ5Yt/mFstwsROk
7GqdY56BRSidgPEKVh2+ef9v+4zK2BdybbA41+33twKD1bEgYV0uJs+3oTWMLezQ
Lplv8XPHCNSWy9MBkSE7UXWxIymZ7YVmSv9HfPIQcBPXilM7pfIdPvSkbRRqmE3E
fQdVpVhOrnFLmDXy6o/g5LuhewHH7MRnqgQD5G52QYKsIhvX2YERWDn4y7LxscsF
nw87gJ6rPmr1dirI89TNsFBplnVxuHIDuSwOgXEyykBMHbXZQ49MnIqPLUjzrQNv
qx4Zutvcxs3LT2NCSA67AfluHoYv84skJwuemwAM0bu0E9h0sdklS3rLLeFkiWnW
LW12anTaN6Xgkn+b/S+OR0l1qDei0tLHr0va5qROnbMbRI09Y4uzIoIVk5RZk+D7
7r6+UFeZeVUQY5DVMpPY4s1EbVAsy7uil7/m4iDl23tKgq9TbBuyTM7tCM4639Ug
rcx/ADym8IBRlx3Q3JKmQy1stz95fA/lMEr93u/+gpYv5SLcoXoLK5hrFaibfs+I
3NMp9jI+zeMz+vODV0s9E1lSrI8YHZig6bPRnL9qQ6Jj6jcODuTqcGVtBBJ9FUiG
raryqngGf3/iJhyWl5RyU/96GJwqHvJmBhAOws49N0zUXAFwhDW5IxY8u/qQQgS3
3wj2NuNNYB/2D3LyXZyiGc7ngi/osHBDtIWppi0YgXpWKOSIQnVnOxivdk1sIM+k
SaMcAopjtxYsrxOJ7G+qTQN5+c7mVS4DvCLGNch9kMMb0MUpXJ90q/FhD/Ept6fU
aVdqdj/xRTWCixKEPNEcrocA+881nHzui999BsJ/XP6vWVMTIdAddCZx2oZ5Ca12
5cN2yH/9w+vO9Q6Vk53+5UnroEkd8y7z6zPGvYDQ2EA/31MM63XzaPkQYPXBjZbf
D4wGYdc8vtgl8T+pBljJGUH7RQEEJHtWGO79BnnBPBaSVE1coo8ZzUGY34m/jz+7
uA2VBA+aVvbsIVsvdtCbYMqK1y+Eb4SyBg8Rua2F/HoDSQK7LgTG6eOWR9tNFU57
H50+05K0/GEe2WNrg45dNgyuBgCbFqhegd8OJPUiIQnHPSaC5oxYqiOMxFEXCp1+
GJYpCfSEbMi3b1+Rfr4ZvprED3oo790E6oNaofDaVXOhUML3RNosVZbb9y0O4rNi
PTHBZrvSKltcdnaC0M0bnVzrRs0EEOGbccLu8uIYKRVxA7aE9kwaRN6PcsIP/WPN
QYrJD7CgckFxiojY9z0pUxQZVJw4l7WSEvKc6FsoQxRUNIr+yh090RrPI/XExB8G
6KeoPpW3WFFUjxx2caM/MeJ/UxHCbRIaT9HFswK4W+BE02152DuaIt3TdlHkSA0N
wztRL3Wm4jViG4iuL3OeWnzU837osByI3O403teRSCUCqXmiHwv9DYGm9lVbjnXF
bIjihLF689nNhvEHwsCsx3Pc7JnRqJRzEsl/VNT23qwyP3TpBVK8Z/AYVieqGF/P
cr9ehYrcFVJFkBWZWE8Yq8ABjd9zyOeR8N6QpXfCReQNdwmNW1GDuAxyqZvZwbHq
gzS6SLpLwaWAkh95WB2egQdmlaguRDbw9C98SF71r+bgwuochGN6YG8hEXI9XWpE
0ew5sWKFAhk2BRzngXoB7516bCMVJDttTgVoxBSGp38g82XJ6A4lIZkAgqaBGYlk
DmgrA7Nr0doznnndVKpd6Gp5v+WViQD3hPH8UFhFTrw2NERr8Pg0wMbfnh5yHE+U
eHTyft0unKl/Z8nVOnEiWiiF9H5X9meTs8jUKDm5znrWoH1PKn1yn1e5Z8hkZzve
5sLAvylZgD3Ag3wmefkKYGXwuSj6j/YOzB7oSNoEJNs+MT9AY+5+j/xGHbl/5zu8
OTSsYCGI2AAEXom3D+x0QiOGh/mOS55dzM4yykThmZLluSp15j5mhfPFcoRWt5k7
fBfvqo7DbBWAmkzqk0U0+pUx1zvNrlV3n4xjMG0/bySsnwGuFuLrCSvJvwtHEEqp
vmE8hRtejqAvJgfH0CIUl48/Dahc8uliixSSje11dF9I7NvxL/dCegMFv5FRjgBy
/m4CP8yujpYg8EF39MbpSP1vbWC9JWdVAmdiaowgani6DvnywMaLVXVbXZUhrqv8
SmVGXl3njX/2AZUu+KX0zL/XqLN2THfk5/VXKQmrP2+bQdhrlfm/l7H2NiMiIJm4
MQTY7WpAj1O5cN/HEub8wgyjpRtafBPygaczyTUBP5pBj2P9LKYU8K79aWaPKc9O
ureDsV0lSFU6TTfBzFUDeIlo83g0e/nuCkJiRK1UqH9ls4tqkbJfqnp5aknsW+16
+hQVi4e5usOeTyqzPHk4G+NnIphGxvyv89uqiVe49jhzSsAST38e7U9pqsKQYeww
x/IjUD5W+ukU0le6rTZyrq1bvaMCXkQYUZ505iA60BJ+4YiEC+lOR7Qj1lZzYfEr
DB7BOlpuQmkjNz4KqN3JDdMBrwvz5wozlVNNvILNgVPmvKkS73f+Ei3alm8UrmIb
nn040CI5Vzko/n4uBUBLs1RaHMkocRY41BSvgBjR/pGNr9JJto6uZCX4cbH7rsVl
TDbgw4/rWwqeP02oH2XD0oLjymaLOhEYlMPQ756KMk3LPIhNZ9kvG4TUvUIQHVl6
D2x9WfQRNBIrbSon63zUvhPLNDdHeM5FHzfYlm/WuxWex4FNML+L40ipZX4zKj2z
Ze/tpFlREjj47z4+PLKiLzVaQlkWWG/+kPN5C+me1/UK1lxs/gtbyEAdlgNTs8tA
gBaneswgsCgvkoeBJhc8GgWCdWb1RnKhyMFFQNu0owjPpTR8vsrsbkkTm6sLb2bc
VbCTWD+d32zelb2ufLd0oGmzQZCh5x/IhicHUPT01eM7mWtbgDt91KiBtW+GfIwn
/XassWX+CDYarsB3oADmrlKyKYCFplPgDgHHZgItvdQtlfwU7Qu9XMj3EEdlVjcC
GgeZ76ai/twfmEqVRVgzB/DXbtFFVfiX7g0dUuDX+mSm74GcDmOUmuslHZ38ZEF7
p7gU5bOXEFcsGrYhTm6/xMSXDFb2eLoyX26Rji8b18EtSeXkCZhRdSF0x+QPi5Kw
cRnR4dwyajpoiirr9PfYwLuaBNWN59gYFQiQpFVBG4iAVs53hktjG82BYQre0VMA
jAgK1MCfxuz3CILUsDO7yGfGTXtqqsLPrlOgsTQ0i+0FunJrcN2hHJGMLp8zdrwu
yF7ywguk7o+EEd/T70LPRmAJuFzNkRptDTE++hteyx9CUJM+1lz/uCeGZBREs96Z
rkC571AIZeR//Ka+Lzco59sZ/zyAGe4OXrMV/4juYrcSEDrglvpl3NmcvXquBgXH
rLmGsOqlYJplwRli2mbcjDWkGoTwR55szcuAEaGydZNeA6UGYqX2uJzEBTZAUn9y
3O08pstqs7/pXqNKQnOUpEfPHcJiknuzrV6j2XlYr+R81apVY1AFQRpn5JFGUcf7
hHZxXEManNGB87YCmhTFYaeKh2tVO9un5ZzmgBV7ebOtyfiZ9m1fi2fgodwb2iYM
aw7bSzvys8XFnktKA3n8wkqalyEkKmK/0Cg+YNbUGiU1e077FaFs11eFnxc1gOOV
3Dh8RREygorpHvKL0Vep9om7LoSwC5vg8sHxeDzMRq0AaA3hyXnK+/ytQjG8xzie
Xehr1ETNK2tORwH4HKInf5hlAnwTL2LH3E0pjQRK5zhfKKX6lfg3TrrQN9C4e2Fr
1vEbF2R5/MbwBNHiTDGE0sdZTFA1L4i5caL02xWjgZwVLfFtt2ZtccrkZHFtvGZw
9b022pr1jTjPlhkCqXmEK6tDOxXjjzOt1XTYSNGgh0wrG3LJvHW/yo9y7HfQbO/9
PUFjgaNTWLHHbKbDkAeu9t5okT6f94rznIdvF9/ae8skePJJR8RuDHODwUY/79vX
JJhFMJLHmlmObVIaKKnjl8UVfTEJJWxgfqRamymSAW3eSWtCvZEsC2mGjJULbDbB
Ehus96eFevZleW7Zb3tx4btI0rbyfDDqhbCRu3aenud9nd4ybJAHkPdGrgYhx96n
p4qMZAQ47h/APXPsCUQy7shfCJOCoBweB9+zWf/ZRdjNhS0BcUCX+nBuQw/JcHCv
+XUJsx2ySNcILFIB/50/ISwFh8WoDhpAdxKQldUaWt8NRFlh5rG+n5973mjMxUJ3
U1u/6ZDuhTVquIomjk/P1P3rN+awe10br9pBrcm2heddwM59cxRgzDJ8t8DoWis+
XWUfWndckx+bg+NkjceYmLBufe0xHwTKyCXYP4ivZpUkYFBs14aH0seB3hrd0URM
rIwlJCjeEQYFqk0ZuRkr9Qh/XiOqhF9GPjcQ2YO4cMYwHFAuRpfPUsMX8WT3ZVd2
AXx8/9RMum5zx+olhXHuiLpIoDxyfzbkWZP0D+1ZPROlq3n7WHbLHng7tAIuzl9X
UXTgd3CMQKU4495YhRsQ9VtG4dUay+syQFvpzaJRSVhXhql3QjNfNZ4FjnFMOSDF
2H/ptnim1J5MB0OjGFd0L6XQIJw2xNcr4tUQ9v0zgSfMtwkR46AQqeaHbIGgILBG
QOsb8jKSCjgor79qTAqdxABL6ed9NeyienYUOMCs71Mjh0L5oCEX1Wf978xav76W
061PTDJMYhsFZw5uYJAVsISSEX5UGx1UGX+nPMzt54uAETMsbg7b05yzw51V8Lzj
V+vmZSCHwsryubAPwrwqoSq8cpHMOoe/qlk9blbodwgIiyIhydJooPuzUCHxsKFK
o1ahk2j1QvSAs+ubJntHJ4yeQsqFNRrVBiHuZLWiUpCPPHI7mGOMOiJsJKKysuXh
z6Gyz9n1jwXHM0Y/ic99P4uhrKiD6ZKTTZosDJHHP6FescHyWN25/oz1hrALHs7v
uZwEoTO2hwm7qxhBdTsH5kPczyqAtx/JBhUyWZQ7JcgpTZqyc9g9kBc9rq1n3GJ8
s4NpZR4yBjUADMZHaZqWWx7i0Vxt5M3QsIOrCy6aVQpc9r4iu1MCIK6R4eOrs9X4
e8ZkSHSv2BZ+mMbPy88t3tpZ9fwgFagh3vwRQUx8zsX7efiSVP6D95yoQ3L6tgoU
JMprARhUd88wCFwc/XXhJ3NcQ6libG45VGucHUVKyfptRP6xkXEQm7jio85A3xrT
RDbmVQRlXZ2CP7hrGR1oZJSzvytogb4FZ5xSqc1mVC1crsm99jH0PhTBfCBKQzeo
l8UiKdh+YEkjH7bXPUxVeN54PX7YkpZE2XJtnNHIEn8c/0A72L5ParkiMF7wFKFU
jROcb5cRIOYzP+2b5fKKnIpiYLXs72yVvmisQcboapW9AhrP1W+il9nSHhvlFbVu
UFhV5US0CiF4CffCvbZiKecH6642SuaVhaQNohCCu3yqEf41kUoqAZGW65miBVCH
T6WyUqfqV/wv/Cy9Bs7f0QiXoAEe6zXxESYFS0n3LMov3IZi21LlY9FLH6Rzelv0
90nN8TGozLjTJrJLPHl6QpdGB7OQMpHd/wf5eSLr7onHzsQqBc0/8FTZG+WHRIdU
2WfcXH6SBHMXm6WmvLWWkkPXyEfcPDdEXc07V5jxtO+JPRtiSefLr5vQLZtRVoNW
RSjg1AEnikPcpsuVTaDXEL6lhEqX+m/joCh7VFpwkOG8rEM0RWbLV6GtVqPXL+QQ
4Mna9Lznmc6EczRLX0xyhSX1HWAuUewGB+AADocYKNW4yARlHYEAH0DF6WImRfQe
hLbh0QL6ZnnGAeaSGZXFeNxg1cgGq3ZF2Vyu0wmB6CxxLDcSZhXVPsvibm8/CExv
3h7igM9vv7EJOQmOCj42znEfhWkyGnICqW7a0zdh64aUWo//Cdj0duT9DkYSS6U2
YXD0ubOll5NiwFgCgoUdmQavUgiTlpGp5IUFkOQeZY+l6X6SrnUgMYLHPdc6agv4
R01Cs5/f0d8f41rxr7xjLF9npgJqC7lw4xCkNnTheJIYGNLPQUwmVFZ8PaHP/0a2
5r6A/qhGsGcD7PZIGfYfyZFXjs4asmgk+Bzdr3flqfHMRRDsBhi42MVCSDTXo5+k
LinODxMvaGOfJWJWOY9+7FB8LQvHFzH/NYsEI3rTMGt2oqr/lzDmr3RcnXBRfXvs
YgAEtDKe5h0+UookhSOGhWGyogOvG0vyvbRT7V6NlkTMvQtZDIS0v53LYdbcRiS0
KnYStXzOAyLi4A6gFcxSobJrknhtD3ryiUxxzu5D0n01WKXGtEXXVKcr194RkgM6
RfLM3RuUrmeDQqXluh0LBS1OFPaBmCaVUSc0nvOgVfd3wX73R4jEEhCBBGawFLKH
Ap0uY8o7Zz0sjcPfsmq/8Al2RSnd/e4Pt4d5seVOA8BwGjw4Et9n5kCQwvlSgedg
UlJKyoAgrQqMDAZ/UKAK3plcqfdmlRfUeIW2UzYTh3De3OoCCa/DvqP5SgIfi0Ie
UDzQ7hCjgBuE8VbEpompBLLs4T5axqwmNMyLLatvWGqCRjQs1znQ6R7/aAAivvlV
baHIrIHn2uelz4yvdflj30ZV95WXMBXZZExPrbM61fljyIsSdmgu47Xp0CedC4Xn
Bi/f0LxTPDOpLpoowfw7J3mLcfX0SoslWaCxOtaQBkbYNMAOqgTLaQws8xgFCAu4
rYawiMzHdXznjtaEw0+Z4Qs3NuqezQGIOb2sS9Pt/ry+cph2aQDRP1fS1hIuTImC
ThSb87xnYUgdEW7Lv2VNIia9MzCdLPAqMszujtM37msyNy8Zd4oZHSSV1C129gVB
1wVZPDhtMqshUy1ySIlX7Uc6UWLkSryaQb06lkyXIbknzqxyIDbMJgyS1w35U1/j
+LvYoMU4YWLLcff8zhYlFMsTr09wwPghYF/FtULfLTznfpfZ5p0r1avAhTttmSCH
hEOGPHcNpcr3PQKDfr5DV7oSTq/9wquzSFBt+rHG3zDgdoM7+AepY8LN1u6eUIfE
HTquhUQsoz9Hg+uitXbJKckAcYZSgMoPgvWfR+ZiSGh9wb6H2gQg8uJvrl3TKs/M
MHNoNRFumIpz7Wc9cBuCo4Ug3fE04zKx7kB0m0SHD7nu80LrXBh11xz5kJWeenM1
35tLJEzx5s4eyWQw4V2lnncCzsUiLccLfk1vvEEXe9SI0+YEG9ocHpD6ebUyn+B0
gHlk68FYLofRJBWZLBYXJbMwFzxbAdmd57BiqEQWdZKaF9yBky2TH/ufBUwZP+jv
oRGMPPv9y94IiNjTOL4y9mg8eYKQ1S3fOCEJjoby8mC+scbHUhLJ6wcT+YH7UvIk
BFxeU4nWOzqmVQkNHvuCLRlWilk8NA7BBuyL9tIF3WB9YdCA+xLCfUViF0v+CZCE
gVwRUkFjp0XrOW0mvpOqzXsMNvZfbNAUPJjuIDnerGKt3TBpg9NvQG603ZXtkllR
f/u4tbJN8SeLz9w8/JCWavHiazVmpmy7/E2lkhaoFWaM6lTyMU9HbkbeFxcbIszm
1LEsx2GN+T+EeKwJyvvOvq5dxTU6hsg0sA1rL3wYHuwo/U5oEsTRc6vkh9HheTdN
CLFDP7Z7szyv5aEVxpMjgWYVRxW1/zjZqhI3SpDQmo6Trqudh2myLLoQdGALg7qu
l/0lioY9trEnrEPT0bWIlWXfhVWTD4CrZJVbA+xr7o5cNNtqDL4QCbSCAZjQD8zG
XnC7JEIr/yiCWowCI1wwHhL4w2SGM2Wr4h+d+AYpkAVhuNfYPZFwNVF4FtpRr6on
H7No534MYTYpq9uzBUa55OIc+s2I+H2YXXGKmNPsJh7VbZ+h6El1N6+aAthnrj8N
0b9VRRMMOAGsQgiNzTQVY+5kDEOwH7B55Y9MdXMp9hyH67rbc3vOWLtsC/HaCaiV
Gg2Ql6DWSmhQX29DqAaQdyQq5bkdy2T8/inY0fsZLC9Luxyk1vh0+n1Il7NUbWJP
QmbACd+3ba8iTqx8121WIpORO4no9EyuHC7qAZ6SUqPzzRhhG32ObJW0cxeBKOL5
QHPguf1IlHxO8GdYg3M0SsnGeRXTfcsArZrjhPOdVCtKZmjLnTZa+ej2ywEGtveQ
W23CvGUZSEtFAqiSEmW6ZD0IssoWY/tjZy8PPmiD6ND57JKoG7+EIxmJSO5nV3xs
+lojTzhBXYNHWteLr3Gg9v/snpRWAv1JlIv2bo3FAhVgv43DHOYaPtzt4gRE3ZZl
60UDJ14YVFcJcZSw3MB3ZTiZK1VG/vGR7fMkHOuZWfWBJ1TvRbZPeyyvqboAmN/P
7CmnaJCejRslf7eGaZ+1ga/5B+GXuSTlsemBw63MEmglNItQhMqTZM6QOdxbW9lm
/RlM/BGfxTtcBUm67J+wxBP4yidA25vQBTU9q+BYJPS1IdP+KHxCqvYzGXNWd/Dx
3s6P7Akqa4IQE+/URMSCTiyiN0njmudo1VQV4t6JmMFMZwaxO5byd7zjVQsLr0sN
IulQ0SpdqY1w2JkuaC1UnOVtF8nJ448JyWR1hUnDH1k0QZrK6qHAvNIqpV5yvr9C
J7lJVzdhSIj6+dpZ60VBRM+YOR91WCGjCXCEtYvnaRLKRb8pxUq8aT5eLfswqbkC
DglMwTX2tYCEDF86Wph+jUTxMNXTzSjVNtu90tMIrLnp0uiq9MNY0sZAY1ZCt5bm
Nj3DyC0FpTYgzXpHT9Wf8Dcc2KHL92omy+OVyXcLmJ/Mtqzr3t18qZdee6Nn3qsr
KTzzjgDfIIFH5Mn6fnw0H1qiyFPzwJ6JhheiDXi4YCZ3hNr8Af+BsUrU0mAiliGL
ndkN1sNh3VA2ZPXGnMJwwmpKyzSyxadxCjFlBGUXrS8XjkLxyywoRB+s6zqUnu79
lA0kqa1Qi822cHYQZp7+XvuYpZjTY/SwpDg0VHwE+hnjrADTtxrXgbgitEB0eYoN
jiMhcEU6t5SDZg+6rJE861pbRAjKb8KAOhWGdg+IFEbrY6BBXFloNed9gAyq33Up
c0AhdfeZQ5IwNjS1rm8+KyW3qw8Ymq/8yBxNOUSuNKH7V8cPZnmuZdzEiosYv/Q+
V20wT1zTGljbEx6igtQnu7mERMzUYaUKHyUc1NJVWQSpnTb13ZZt72G+Kpj7cp0o
qrpBGqVZ/W92/GYDtnky9xBLOhWZqOSoa9Nvhq4xtVFy8hw7CAXLvGTiGYVECms3
4V4vVcdpS37aYRwqfjLrilxS3DwOf/PKXYl7m3RniXvBdM2yZzrZCdM07laPbgg5
r5zwIU6+P0kx5zeKOATZ5wGxKxYOxiegw+ZbWev9KrpVeogAEBwGicLc0QIbDDMw
MsEL2PM4dsJxNNVmm7G8upFBgKSKFo7zlGX0wpOPzI8iwAdwoKkT3/n7Tm1Nmqn5
GSNlynhbHuCH/YS0zwO8YbttvgyBWB4Li4db/CwM0CmPj0EX8eXUkk82brZjnl2N
wCTxisLYwJ88zKT7rwLGekVFGi4LDutvG7Yfwz0pCUqiHxo6x06LcDmwAm44b2cb
V45HJsfzUpsorIIZGq25O5H2OTKJUmDkn/7wP/eqLxMCOW6Teuo43Aad0HJ5yqll
1I5nX+rmUacYcwRlwXIQzOcPyVrCyWPiuxS13L/xyLgtcsFegMt8Zt+rEmHGstFl
+8OV58ZmNu8QwUoBQRY6We+pA/ayqDLBP640bC61bAlq5tSst8Ud//VTXuDXa7aa
L3ss42kbOTwIb8kcLZn5AUgNkrxFlKv1gWM+8ElmP/2r+kK8B05UqqyUpcaVi08Z
FovAz/N8skTfn9S7RT5MULESoeoozVA1cTFOsrw1NE5aBW0q/cDJnWgDxPJvXv2r
3KNl4qHYTOszxJgUnZxRiTWsXdgnYjUSC7OVhMmB2BYkoLavS9XjPgtzDYaBViZ2
8IyDBnSKvhpg0T+xCIU0EKEQzoGORD7H1jKHNOsujrKfK5XvhyWt4ToG2egKJUQl
7RUePQlZzZ8oWVnFVKaYUX0ngl0x2byXfkFcWNedLvgI4W6AbA+hryjgkK1nYfJp
GGO2zhSYi/IlZWWHB0pkedUePlHm0jPgwGXMvWErrrc/6FZIP/3QJiz/eGGniB7D
RWoSoqlLFol/78HJT8hMz53p2XhEcwaAEEKnJiN2ARuJzcFG/8zm0ILUNsHoXsqA
Jq52UieGXV5wMULt3dEAztqqPeK252/jFYR7OaFnFjKwm0olEd2a8bix2BhuBZDZ
bGyWaRt65MBI1KsqpdW3ZW4W6+1JTuGrlig9BZyYD96k3flKw4yrDV5484njGxzb
wbzZmYfprF0u9mdsk5qjpbK0VoKcTgm7Iq22iwQzv0sq2kv5LeAwZ243Y79Rtv4b
THpySK/4McUTpSDq7J+4zHCvHCxmjDHRclMAxdda7RxBiucA22OcxbttkWAKKYCn
efIsSRzXUNjZq5qT45HUBzN6ohInhkUVlktJNi9FFoSJDoJB7puZO9pSpEnKaCuC
GmsotFkpgU/lxCBw0omFkuc+QAmLOHmq/X8Yo1/QyiUwCCm6ghlEZoFn8pqdzpAx
xdMSYx4sUO1IMMDjZJZSqFDPkfx4z8OeUpXv9RW38UG8qsDz1Te6qXrfDc22rYTK
KIe4grpMPwIXlR3I8/GIYA6e9fP1I1RtBqrFkKuKLEFrdwUz3u5Ux70wprl+dry8
cdSpgjmHrmJL80Xfqkl+AlEQ4C9dhWqTMRhGGLcCaHOkBdY5zy6wX09+bNj6DoMa
CaH/gnVETDOCAoY5krwSavsB774C4Q+sFP8+FhoJLT/UIqxgby3/+tSPPlKT/NyB
gqBgnNJm1hCn9Xs9e5qREseawSiI5E68w7efC/uJHxHytB+oLFBLiKGgz6tiRnaR
bIavLAXCZybnRGXeZI+M962ltjJqYK8YTm5glWT83kNpMKGVQOeXrh7bqXnYhCHM
DJiMDWENBsQlAcIKYusIFdt7ZJWrxlAxggN3a/fm0NuVn/Fyv04nMFPBPR2YoN8q
eNs+erFdbgsoIL2K85h3Z1DSLP+fOSmpl21RpAnNdngTUoWI6w8wqghQX4e91JVc
gQZPJG/ddb5DAvR20ZnyKWNfV4aR2zFqimCzqKjiQVtTa4Ies800QvVsigndlW1y
kSMocu1+pTun5ABvmdkd03yeefoSRQcqRsdF1W8zbMN/lh2sl4Js8kj7mU01Dp7c
n5joawvK/9Jsdb5JR+qnqrrN54scCQ0MaJWOFulJQv/Vs55HlsK9WfRRP/hpRLW+
Th+fL4vVmb7S+Sj9upoY7feZLJT3czqPvWVr1ZMNIPg6OaDZKR25eAYjggagFdDQ
hIJJkEewIp8rvgD3RQZ8CSQwxvuxFsqYzr8lUzLpxvgD4OBxbW4aBOS9K/QUg1Rh
2WRgi4uybUHwBvGOPs5uDSlrlq8G/WFq4LAlLRY61aK3+TbsDo34jsFuCkZOhgUl
AQBZqnEZUPcEt0Woy+gnTvvM9JgiwOWWOYuJc6+Epq499loI7C9VXpiqq6WkLOHm
CZcrRPwUzzAWtxc43ibaFsgk+MJqQkQvUku4Bt4kPVEkHBqJhcRFVVf7r7VHKkSm
ptWTb+Q2vyNuCIecc1IYOPUUZ9yah2kNmvodCX8VJ1BOpFyuP9DI86S/smDaCWNG
4uA0f4ypzzjC2C+LyuBGOkt/ozW+9CCwab3E288d8s08gOApQ6F48Vx1NlsSHCXI
TedOyyrbB9o/FsFlJ5elB80MTQDK7k7SGlXmAsGsw4QRcITd7F+zs4+OA3OlLFDW
rsUD6yqtLtxTgIMv6jn80ojrck26xI7nFrPSv/Q5Q/4r6k+7lGx/hFaNeanFeOGg
xn3sKjrkf6CiGqie4Bj40vxW03JMgnXbEcQE6xig+1hQZ3/F90FfVQnRoS4ZwbE7
OKwJkIKPXY55yu4RreNOXjJ9vY+7TG1LXAM31QuyJ9wgRgnt1vN1HvTv5xvNIbfq
eKE6FRqIbjyPfwjEjNUxNPsNKqCV511Ni31Hkt54dPkIaZzpmoDMJOdKwsO5PE+T
/gs8XNmA3P9E3JzImk/J5zQ5K/9P3nU7JOPxRaZw1uDFWdLhWoDWvGSnFlduMWea
VsBNmW8KBjgRzBbttUc3X55QI2E9KILyG8lfDsYaBQLNnZMvRy7t9n0vjFuTbgnw
XrlTRshUyCqh9R6WpMO59ecVe/b0fYfQ/zAfTyCq6Tsq19nYTd6k6pX5WV6AwU8B
ua+JS0E0WoNgitqGeq0zFO4+QeuRJToMFrQA3t9qnZQEJRSH3Bqs8sVK1WiGK88Q
6FzCxfdHuSVoZVDQkyybUAo31FbIGMN8Jo56cUuTkEa4xo2vk4KyL2c94IuUdGab
vhlgg+gzhZoxsA+bI2ZVnfCYIOLDNQwHLadWwpATw6qpJMOVtUGOBD/h1i3VVkhB
9wL2K9m2UivzW9UTja85gFszeVuviZL1Ek7ooxd9qSyHxR+dpTO3ZPj1vfokfNlL
fgMJziE8Msom+ug+L1QjtJJEDqrNxqfobSoO6LCyQDIYDcBFOmdf0ocAxTjhxjry
KgshjNCdVIhP1W+MagmPaj+W/DoPbWUw5nXeX5cCUGNjdVEaL3AXluX28c6QLJmN
7Qhji90orJHhGPJ3/g/g0sfzgmVXBUqUFiNi8lTkdj3i3/j3gsEZRig1PqxK4ws7
0Jq/gcNDjPjEBo9OBuFvfPsGzY1/SAyJvU+VWIXbDKG+B+PXu1J3lDcIwuoNtgWq
oIE2OkyxumGb1E1ZjlPur7m+CaZfGYVoRx0eRUu8tUAFvHZZzHpr3K8jkUpOjJsy
SWL5vDP396bfQhp2UeVKTKIbTTo4Oa7B5S/FLSEjnYri/cUBizJ5ukqrKkR+DaH/
dmudthyqO5AvBFBWQqcMQmCz/b+jEukzB3a/pGvlYa31ZSqk3f5FC9t6Y3AnSSbJ
AZvdAIKjGhrnMXtZhNwOf0iKdtsEelImOEscPdHY+jiEmWk/Ey2HCVW8pcxylZy8
3L+DmurqyMZtDHMTlBIEEm4Tjpu7oSEz1ExTqKwKzcMrszzz4vJsyHPa7ARXhZEz
kfpYqVt1X7Z1gH7haFGo8qlrQ31HlPHwIDmrybeohM5RnxPh0EfHhwe1sJgpJmQo
cjSqWZtbp5k2r+R1qRfyFlxEk0RJN3gr3B/gORcUX5yhm0TfAK+st2uQSjBsnJja
JzAgEWjsOGPnlvqqvB7PZor0I3R6xAWShpKJOxVm1ayB1/caaNa4Rnd4DqibUH6b
HvaKtuSKPVkCW3j2UyZIiYZ4C3kLt3/f+9VQXVEuiX3Y+WieP21FO6X49meqkSp8
kMVf0PoKRGcc50elbcMfnK4MvHoIGv6NzoVYzXh3ZcApv4oSB2eIUgCWaJ1iBm7c
QmKXRv2deBZe1PmxCUuMecXYdnvxc+0+5k1zt8GvkkqAfARiv1EehPSYEJnk5cAA
WNcVJv/n/PflrtsWiacXbHEg3LOT4Oj1ae3cvhHlt3bmELF44LqZ2EcBZ9wk1DYp
O3MVkuua6CBrKEIYmjOQlBJNDR7ceo74qsKMz2glt4w+ciGO9QHosRN/U17wWrJ/
OnhYuyeStoNp6sEsb3hBFubgZyQyoV9J8ls7YsAxbGvKqc3+0WNIJLg9uCzlWRVJ
kfA2dXeShmHy3y8v+iVmGVGjOtYjnCEDmKm0OgIbdkwPVE+/Yq31iHrnpG8i4w5q
4vB+N/1GF64Bjdkwlr8hqhPv7IKKIWbTLJkixq/EjAERKtuVJ46yjB/0oSaXawsx
0EnTYfZHldK+uYQYvg1sWml1t1pxHZkwdei3RaxW3MxAvzat3VSibxWYXyGhO5UZ
AYWOr1EWPbnM4pQMxfL1957SzxxViFptWyQeUpEfAr9ulrtFGey0FTXW8vF+nDHk
WdDGaL35B2UdiRgHjhgjkO/xrF+fvMm8KJhdkI3tRYHabrhdgza+q/nsTnIaXP+4
KGStaAS0uX2Z+7q/IFiiUbXe6jN2rwf2nBvy0y2RKEyFmU8V81H5ADZX5sRP53cE
2gsV2VsfWDoyn9blsbmVgRpuCeX+lLzeLF9gC+DEOpsoTFoDpZL7fY2V7ZgA22jl
mhYKAnIz1TXsL2CJFzAvlRQvDven/bLb/JbjC3dZQnpNyyZa+dhuo+xgFbY95YR1
yqChxQaFSFXhahNq7OMKNaaEzYmNKlKCHylPoQUEc3gJqGtoCXGuQ1GW36V/Gq91
pR2njw0M9as5e434VSU8lcyuWbWvYryDpwUXek8yWnz+K+zA07QqlWGmbjYt69ep
LedxFGfTwJ/dSWlirEWyMuLDzJsdC32ROyKNV0QBRrzRCMyfZUGjALeU36ImHNA1
lS5ihVWqjyX6N/YuMtGt69/Kf52vaHSETaqw1vpH4eRtGx0BKhRGSgU44PU9tRJA
KTrr80UMLaF/7FuHtbfcj2+aTZw/TqCHnc/tUQLe9gK9QcSZJt1JsAVDf5BNWL6v
dt0evL7318rvMHVORE4ADakaz/CJtetjXD272InJ+6wI+CFADl0sso6O5Qu6BYug
AcRgowrXRj2Ks7mZsbtk7/IrDvCAORp25mtYRpR/R9xgz0WRtYCwVAagLlEvPJH5
NmnJzuL4gBNAms3ANKNDHFDSZ/A5H+XBCQ4cne1f6fLQ31ZJMEU4mKTa+DsZdB87
Ur1eDgFA2aNUAlTS35hXjlsN+aFYH7W0Zyhtotgn7RghYdTw9HS7BBv7UBQTGMl/
/YoP0eXnxugujSnz6EyFyrUmhFSIOKyX2RPcWdjMZmUQPyC83qTPxFgXki4VlnY1
iI7PTpnKIZjp7kmThEvDjWcQGXj2cq+dfYaG61tAlHpjMPRVh1g7UjDkhF34w0q5
HBP83OR+/OZ9pK5cNJB+3MLeTaDAw8D1eDuBVLWbXNF6YEaZ1UAfgW/mTvMB8GXi
Vl84h2TOSuaxrxJs8x50ckSf2leFv4+y6Flco+x4BP5kYSY5osIDZ6peVjt4NP9k
OWm34cysUoo+jXCD67Ji2gq0J8zcvQrrA0uHDQcaW9A1HCxiaPi+rwNL6/c7s77K
TbMn/e81d3s+BSydTvhfKH78bFsUxLqWiSg9EXnHtZhRlaET3ssfq3z2K+naqyOG
KCJY5u8Sc4G+w7zpDPpsfv+V0EXiSx7x8SkAP9Hm8yUs3Q6TfQ8XlHOg6Oa4/Y8D
CtM34ICVEHkdAhp5CgB98scPpv2hJgEeaZe3nwXEW4doF1FiSNRYcnj0fVfpbFYR
mkYNBDLz6DYrEUqOojYXXuWcPMt5IT/1/NRqNi3DKwnL3ZQKc4xQ/zClZkIiJpG0
01xYbZeJ1cc/kqfKL4+db12s35//GgRnYhe9ksJ6hiGiMnaAWXUXVOMx84yCCgtW
MhkPa4oMkmheOESCTIKH5bihOfLw3si1V2DvTz7pS2/py+GxZIDBmD+lZwdROKs+
b1yyCsyCn8/S6MlwpMHS7bVIP1dr6LpkNwFvg4sc4/NzvZK1YC3WeBgKSLimprVt
BkSjn57YeSdleoS++nJhKPWK2ExAWQ2+Z1Oi0Zi0Hgq/1RpWe240dlnJUzb/R63O
hD5Dob46xf7XwzIJn/f8n39130VG7khGuzZxhKbnRavXEnUz/GRuDDA2OgkWngYV
U7hvMnSoWQleCc5fkDKdf9X2GLbTUahY6hWA5nnBkdNTH/NSGePE6THZYqd/zdGy
4RlAAIUBkFBYU11kskuPsI8R5f4MfCEFv+AaCzT6+4GvPyS+6YQBqPcohvNrRwpV
835tP1vts2/4bRmeXTqUkDdKqLsMi/1s3MGwk5UpnmiloSmNNi/M/q+iNFW2M8lM
MKmYP/V2ADVAsBNhRDZWMdG3TO7qUDZ39VW3m4LVIj3XfWMih/AOsvHT2rKfg3rH
NWjmaGfFKzILeSV548udZw11eyzX78VkAE83AGnXD4dChwzQrdDxZ5xDPcS1rWgG
Aa9GArNE5RgdRB0QapdmW5nn6E+7ayoePf5Lin3W72WyJvKHORmaULbwZMZ9a/NV
iMRJ49dMYwA/n5dtW16Xw0pSJsJirms44SFzvt+iD2hYVeYiirUBlzy05bhatwAI
2JIG3jVRAcSHVTj2Sf32zPi3L6UCBdp7o78t0pGrnVR/tHm47eCh4+rhQEA+mUqF
rczz+pH1bbT9WacO79xbjJmm1Id8RsykXft/hHLRpj8Fl7xnjUBcSaM8cMnFSYgF
7cQlJSuR8aV1t6fZv0/NAU5MAsAJ/m9QZG0x3pXgwaWUMQTrHXrgUlMiiE7RTm9G
+wP89kotme/Jx+zokM5pNsOJUiYFYqGuHx5iR65A7Pm7FFnEjV1N+CR6yt0nIwxF
zrTUX8z1lHB2LgTIX8sfbQJ0ixCCovKLF2EcApf0G/0fZ+/3QRDS71FfwtarZpdl
l9z7D+DAfaF9fTJatxDVGQrt9UZMR6M8DuGwvYvNrtETQkpK05VzCmlr/h5rLLEM
ChWDL84vEVr0U8zNwcFKoYeTfJaSjOBfgkKiyAx+9jSFHdcJBabz+ctLPMfRd60u
y/RcxjJ867hRV7nYfIhLc/1ra+iFeG7ZpsZlWZ/hghqMc8I8hlU5yLyuo/1TW8ne
LXOO6RKQsFAnGMasvvGjuTd77RubHCxtMM+Sw8LX8ab4HkXHPRvm0sMy8fNFBluS
+vHGX0L8wJq8bk/XbeyT1x6POqKvjJzNQac5FgANPQ1ztMmqj1JXnRYD0WsRRl3B
myhsi+0FNhzUbyBqLhKi8BowWwMYDjxnDHUpblyWg/TFAbC+FQOxVgbag3hCas2O
pLYsSvpyBYnDfRppB2wCC8iaDKGWxDe3lM4/7BI+0OTeK+imNiN/uxXbMSxFiuvL
XRpEvoPHjoDsghGQC4VDYFDh6le4bS30izVmyFPFwx6IBFO5yBs9HVlMbpBbaVst
ygE4IdyUT48iTQ/LctcfRpXgyeSWP4lri0kWg0Pg5o+FAqUz/QFYQo9+uFQzMQEL
1oJD9jMUGTqMoLb23bsVDtMDbUEInFR68Q5qMNYWvcLPTXSEcOurWgAjJb5rWHZQ
0l7gbjRZtN3ODgPjmvBDu0LhO5z7g9qNZDZT5eWTkTz2sorSX3tQ6uZnVOdOY3iK
4dmvZ0pNU4y/cc5Ufh3GhbVjimviy16IwiJNUuwl5hTn/4CEmUQJgD4ej2jqlRzI
aSDEaybNeecxeg/9lJ/UwW9YkSnlVll73ZhfkAnJY5egl25Yc8IzFO2QP4jrnf7A
6ewWGlQEYt0si8MATCj/1SoZK3QUYrnhhRCqFIVWutzdbAZNOD0/bcn/KXQvI0t2
h8qSj8w4MJdpYMhqE6U53V2DmFVvUd3I8eUn2fwPaHkYc5sfIAJ6z5LeX7JPbiDE
8zE8k0dLGoHekXn+QhD5qcafcgNJlMFKKVH9yHzztR2YMcRvZxei8xflFKB/y/Fk
NkSyL8cek4wWWOMQR6V03Qgvklr/kLr+do25x4zZYoHTBcLLVbdWU/cNgG0E2E1k
KaF3agPM71v7eba5uPWkpG0ymcMnZ1PWMRKkL+VsslxwRvPlo//i8+Y6k7tGqEwT
3bPgjtm0lHXKM57GRQ1/s0trQ87bCvX9bUutGEfboWjPRMZLaRAmYLO4g5d+Pvwb
tYNcHmWsTDkIWpFMdAJXUcy2XyIihLuHYP2s+qjiYve2FWNwqQNVZu9M+6hi96JB
A7I/tixYumthtJl+v3NACHVdBKw28YDlAvgjxIzkX4hH2peOEqJdgfPjZX7Saact
AsF6kr2PUnb8f+zX9RNwS+5ufG0j1Da32SBO5ORBzuyLXF5/+Te8q6kwCvZlQcDO
5e4S/WyngQFR8ly6Lm9p4EzQDz4ZY8lO5wsZMtj6QHy7AZwoB90TW+IdLqMz3z6F
Btbas+MzrdeN/HmMvli00F+80ew9YRvRCs7vNkW8nWNsQvYEh47vBeVv7aLht0Ny
ZEoTqdu4jcE04FoJH1j2F8WEUaby+oBvBjZbvgdkDsudET1C3j/3G/ohlTFttdQc
kosT0hFdF79N7mM6x7eoOfeEt2hX/B3IfrziK/HTUiMNKOCwpA9JdTbGtgK42SFC
KIVBa0hjAW9h3aUccSBqGfsExYC7ui8g/9znD/FGnkFRpDERseksreygkzd4EI0D
OW781tuPqxgEg7r4JJ2msOD6+OBlc+jsQ9pruzUJFz75f2XE2nruxCFwThbxpkeP
mDyIUswp8qnrElul/eBFNKuSohAuLOe0JccTdTMtYhrrz3YNMefXGoW3o82Yk9s9
eeTOyiXQYYMM3XQw4R+PRQDUGZH6gGAXauwC7Dn6rBHzSVoBq90Bl+OziqF4/YTt
4e8FtJhO92VNN3wFBFYHtmF9IoClDlXCVxDLAKdMXyXKgtdt7HW3AImeWzHmXpqK
ymg/QRZNsdpqfbIqvE2H4j/HNaPZNzKtmvcDM9Jmms4yO3HKxrOaTd9WUuKI4ZNq
3QvOFqhDnxdYVZI6u6tB5us4gxKQ0WCDQyffHR82qJMM/wz58cWv+4ePel/5sHbf
0Pn47Tn22hBSv/hnwiWQ+idlFHFwoduFvzcLSwsWGlyRMomLcP9oPf/Lr/ShusMg
9zwxiKthdvH4TkZVy2xHAUrpwaNoP+08OeoCQi3Yqy4uS/vKAHiiYSzxY0GuIwuT
r1PhxXLVmM/jizXrDTZ0XLJmHEB31NfQay4Sn4OumjyV38SrYaOYk6rwDFq/j5Fj
9A2ptKryXKmIeP3koK+SwCrZtmVdnm1xckIUuHDmgF9xIXzZ3HNit03cOZJiKFpk
yxSaWAUMHebJvrKM++kIcuAKmNBdh+gPAiU4XEwKC5fgpxYj2VR9i1kUD6Bau3jn
b3rV4t1tOsjAy//N8eC1yJkNKyJPUsynm1MSlbqjk5IK3BzsFvDsuAZoItLtVEmL
Y+XhYYMeaXz/2X/VMz8H/3aXVITN2EWg081SYiWBff+Kc6uxsUqsPW2OYFazXAeg
dqLiveH13Vva89OYKESY3tSNkwh61VghnX5exDZa+6LNtiuFYrooZXSXS8Qi2aoP
Cjc5hHd0tbenfCOUc5YdqnJFIhnEJCgsFWwjJrUqm4BInb0M65+rNzEyOJNo4xw/
pvhDsTvoSo25z8tF4hjc1m7U86cKSAHeGYAfbScaDKMpbiHwkEnx5altJrqLRlRd
1uvTEchzCqEUWcOd18ioWA8eGtWJqTFoS+rYiWvPF9tJMTDRg5VZHj/qDuPUVYyQ
W+JDupBmEJ0Tst/+Pg/8yOzLiqPxJlmcTAmCkJRtM1DxWz6qCGc+ypDsL6LEJAhv
V4X11R13a6Xm2DXybmOZP10qXA79ZBV3UP4eYg25hWrdnvGAO7rr8gLZYVSnYoes
7L7PgV611Q4WBhhEwqQGdDqqpiRCp3AkkEsNl5tZ+rKQc4OssCX0LXf7rI1wROJr
gyIqZxcBAmnsmRHuD6N92WyqOsQhCVi+WoYdX6fgij0fQoetqX+T+FdoMAVqHdEh
CCc4u8CD4D5bys7DidrL8sYtyLJsELpynUeQyhNJNKgGzGS4sGcp9aJ94ywZ4Tlm
Awk09o8wsX8IpDt1u7+Bm3A/ecAVenlv7gNC6NdVyaDd0pyYGU3x8ivpq4Y9FlUg
0wBHI0FjtfgKZlRJciG6g9bOP4M0s7tjUYL5ntMGvvosFTa0zgUt+KRbkQfpSHiv
9BGscAe+o3nmlHB1wv5EmKkbGedJZrQoacOkoUXtL776mowm4Iqvo5MyR6a4to7j
TnjmFzK+2lb64ot0mmcVrhPBtcZfDDtDDaZUhRm6Lm3NFlw8bjT7UtUfM05QHg7r
NuDZxQmm6wXG8YNnX6Idqfwr+5StJgGmiA8wFELRlj63YLFdClomkadPdsqLDqNf
oo59LltfMUqh4DRLSacueuAwweU10n6S6HkOcAkZ1MwM43sPF5ya8Wjz4kQazc4s
BeQ3zUbRwCb2Dg9+aC6Zv38rKQ7fQE5g5AjEbTtMpj7YIQH4YV9Im3lAk8c7xZJl
FYw+8YtWG85Pygr9mJX/cGaXXdpFceMBfISUUquW/IEPqnPzqjfO+M9lnrkF+RoL
tvb35do9k/Dl+SADb5YW2Z4djrI4Pw6yi5XX+oFiBoEbpHfbtFH/597zOvtwbSyL
ssPtYtn4GKu4TngReNySOI1TfBrmV2BGCrLsJUAwrbMQDs/y5U4yTgcBRr2gaEaI
Ef7lc5pprwDNaGc9EhcNi4BybICnJFCRlIUU8ASpvieTKnai8pipDyzMHla+I2/a
ZW3AjOp1s9AFArIL+YQ0ed0OdvKnYa2nMJXhdn9cg/y3PndiKiGbh+vg1cRFRk8J
gB5VmZad4NCY1sW1vblUeLre9kLbwBqvv676B4kem6hBQQMcz2GgGVTwwfVUuGZd
2Uid7pHRmNcYQLwCj+AwnBI4hR2yhvTfq8zKsQyuO/m4iT0tubcoMfoFH0GCPUUx
SrfERVELuHjFGjyjPsP2hzwIjsQqgd3jb+Up3qqNOTBpeyKwXatt4qAPMbVnb71i
w/29LgEoRvACX6AUqJjczNw46XJ0S9eV4/P48L997Zz7Rq0Q2oMVjDyMKnGZ8zIc
+7ND+qgOMHdBu/M8j3yZMrrjskzbAzjV91lt/wXC/NignU8EBLtQaTroX98ucUG5
E2Hm17MHXqT02ja+SpFUdfW6A8RrocK/Rh3wXqeMei6zjBomMUilS6Y80Mwwuf6I
DXZpTUQi5itVHDLTELXbeSO14w1TZ046ZFsK+jJonjKiqg1M3tBgcdy9U5Uv0e4Q
jsbxs4HjbWcb0Cm9bhYiX3kRjkn2Lxg31xjOi12whAOSrp5o0FbIuDzjrLT7JesG
rXJmHyl0WdJAYQu9E3ZSsqL3nR5M7ez7TZxiqsdB91/gcbYbMmCLYCIZ/7vwxE6D
F47TNoBP/6OYSrG/f4k9lUv4s1eg0pkVF7/JeJWRcVMFH/HXGQXaLJUFAHUqVHhB
bGmfv+OzSSew4MzJK5j3kP+HGL3oq+wQ16jsMCI2MO+aa4wDShtqVPDmCKaaXI62
4sBzKI09TVnhcIJKR/yfiBeF+240KOELLXrvj87t2Wwach1lY/TBERsZyVmN7a4y
58r4Ib5NX4YKXBTOL0IHsUSHfdicqVtglqkbMiWy3LwCj4rpCAuKLCGxY5/aZed/
Y/kr/0Bb0DF0nuVWt88XIpSFx4KpBiMQMxWK2irTke8hAjRxsW605KCxnqdEotVR
g85uLpcrnUxxRKNlw67LX3dwecsK1lmyngnYFXQAMp4PXmj+12xPBdhOUSDJTDgR
y8G6Je5VktLVbjVWVMuTjNQTb1lv7qmb5pvhjp0mfqoKz12n7jv+EHlqxzADLuFz
h8nzSrrJZjeH3Qp0tpdoAbohFOaFXafaMg6Wn+MaQ1KZzi5dChMa5rNsx9c7tz0G
D1pyw2998AGqOxm+b5Ft3OEvjnJ/Y0S9mPVBxRyOJnMugZAac7ugk/JnZH27Lo//
NWJjyo+LcWdLJPWtn8bFaEE9bAzHrYcSftdYDiEz9LL/0TmTmnATPSkvixhcLyrR
NpkAU2MJU0OxZODuJORnFd2DjkpmZ40toc+6PbHi1rnBip43wjNOMv95iHimbhDE
3ZkI8fU+fKwqWsxidj9Sr1fzzEvzb/o7hxHhX9O4wht2/Hkr58R2dyWCvGzLXAZx
9+0DRlDboGuHEOSifCBvQ6j6tMjbJBK9TTOJ8sd+OzNN5K/Ngt6ufsIVx0wdsKlT
U7+NyuE5V20z0ShnXIecLF92+8mPjwcTDpNwkQbkO5dAES9UsYZ5OUxYUTAzC3Az
9YFFrVBCrwauFNYN1yVq7n8IgtOr2Q883/vXTZeb/NRdYEIHvoT8oUC4uYRg4VDA
IVeOEdcuJ+BoA4xcQrEDsc/RksmMB5UATT/Qpn8JgW5h+vrXIlw6aMQ2nS1xT/Tp
pMNULgG9aYihQTfA2YscLz4TlzkEw5nun1Zfn0yAjtQwa7jhqAb3f0pphnw2ikVK
q7XEl0OlBy+UH6ytkxzybWLeN/t7VjjbZddjIeRn0KcmgBuYWiG/OKj/wqlJj3v5
quDMdJ8+j7g7ShWHNMQA2QRXM6YJQGjioWtpi8XuEilWVHkMzWkAe7LEXE8fyLeM
dZy8AJ7yWRl8UH+pXHhMLZOvctDBkhIxqDJ6zZddE2sTV38bCNjb27qTpxtf7RsP
0/6cT8L59tCGUNEG573Sp2TFaVDn7BGjCt2ef96CCslpcSy/UMNQPl9XQmvB/665
dX6vaJpbKjaTV1F0ihhONYp1g12CkjNMFGoFo6xHPLgr2LzUnNePlxqzODtkwjwz
KZc7rJQG62mZn4PH3Rhik9chINn4d8d1JJT5+jOd+Rj0vxZk+wrjg5EQlu/QutlR
dsxZCfNlHhotG2UQ9WjcViK7sqvF39cqWPnyfPwRo/1I9bsRHZLeRJHJgyUbMVJn
bpY9hYc0dQIfvQIy6j9o2hiSkONuKJT5SJSrVSF7WUruJOXHX11iRPT5GoBrM4u0
ZyaWXHy+fnCDsiAXROF3tRU2Mszz7pmUnTV2UEWuejZADcrUvF0P6g4G8BgNnNdZ
tySZ1BvXJkGrJvDITVoKkAR4S0c8L44OOyXySIZaeLDI2ly2mIg7sTMhgheG9hIA
pu5/KMxgkvR/zPbNvIr0KyOoIAHsdQLf1OJcigP+ULHMgPabvzYruKcMVaX6o6pA
Z4ke42Kh2drwvf2CUYb/51TGvsKzhN9ixwdgSd5Z/2mrvAqNgXYkmca5n+fSx1UF
RpTNHBGRM/2NeDohTt+j9y9WMcijgU0TX15jF0PZprp+dKnE6Ut0E+ewMdHGy2V6
28qFKyJUSpBRhAS4uNL8kR9lCL+xZ7Iv53sx/HkKS2NVjbfbYLvfsofjmoGSI5IZ
sUMv+FxMksdOg+97Or5sJCEJyviefAlYwUtdUyloLOueLinsc29kR/vEggk3IN7P
EcRGtWonCEaVKf1vBtaUMWK9tfXE+pPRfktHOXyi4wYRxBsripPLOKo35HNiTPZF
uxr/tdW7Otkq3a+HCt6t/U3cc85g2xQsuydoS4ItnKb3vHKNThILSQXZSPVkjdkK
EySBVagZbXIzhPX9/PZtF3BFY4me7VJ2pmF/M22nYVT0ZyiXAheWUpy8yKQcTzXr
VCuQ0vSs9O2t62sIEC9vXV7tqG3boELaLUA1In4UvTZ/xsnYKKs0RUYgWDsCn5Pr
Zxn7xut7kMwb24YhQbV+JysGXUmgufNA+2Si/t3iWa273Nz+AGiv8tAvP2gxm4dP
pojRv7w/HBYxw5SQI2wAQBIVwGcMGU88AHjZ/61f1E2apeAduzZlPOlUWBSeKG2h
63Vv/u4z6DvHaoi7OvRdf5Ij52M3WXzJPvA+6sd40tBsVk6yASrlc9G7T4/rk7Y5
5iKFeLzzbfaDFqlo8fQ25O/aUVPZJKNedC93h71f2/fPjPY4V2r7TM5UN4MXUAuw
M/IH/WHOC2l3KCCBkqS8nT5I4fMp95iA/Vqii2wYad32PvP+zCCXBFW0vCQYcCnC
FmxlpbCoaOm2WyqAR/EL3IbcNf7A4PLWAgeIgdGQmSvPiewJM75TOCfdQQ8h6ryS
4Q+C3nGpeOSVDkCo+ixVRnDefpNaHzjPFTTnSj9U+0h7SaP1zH2kWMkHOowAyCDV
f/iISVjE9hXmNe2Pa6kvoOW7ztCYGtnNDXYlGXb8gPvW7sOIZGbBHmtyryu+7JN5
RdINPRY2O99jCk0OhVb76rx2UzWiRmLuWRNxiiogsFsSB0DHN7OJID8SbX6S1/Oc
K5npY32ra2gnWBDN9hPeG2rCsv+W7Aj5mlYRzqHBkY3EjKrpKtLu4+NYm0ohH3Sg
llY5buNNzvFFgJC0WZd3Llb+Ds4k7z6HL80XJ+DRI0O6K/ls43tyjHjKGrYqpYM8
kCovbwqt+sUjtEKc2IVoSnCKGDwFf/9MH5PPScmkFRFhRk7f+JZrRJbUB4/NQvKF
ca0xZF2XPrxljGhjKpNhMyfkJJHm3f4s2TjUkLe85cBZSYDzYnL6s2a+MNUDnIy2
HxzrMGWY3cg4yATCtk+3nXH0ifhHrtUYlg0t/SG3aG0erOad43BTCFwJVCjP3bXP
V9nFbdKej6YNRfGCIqH9J7uFJZ1dPPufkREGDTlatqOj2riEfPiJBimghfeQADr/
qp3I+cXKaF8LMixqh5anZ3TOtx4smPeQgw8dvCopVpDJa8cryOY02fgHZB+xHatm
UEbfCoB/ln4rtSVQGP8SH06PDdP/J6V13irzFX/qzji8BMVq3flJI3v9bkOeMp+U
rxtb24p/4XHpxPkqcaRP3dhaTvom2gFVtTey9ZY7r9SAaFd8jzgClzIP9clxIAK/
G6lK3d3HU1b8thnE0CoIOnqkgrXOgqMMy0vlMKXHZknOmOM2PxAY8qYmP/rp0cbz
iIB4kExCbJZ+EFDicTDW3Z1L7Ru1uD+9gxPAtWuH/r+MEW02NsB51izEeOsVN9iS
FpJPWSkJdcZgfNxZWCMcg/EaJKbs5L6Bgk7RAPZ56KMxSTaUDe/0D6hK6H5RaDnw
VtiNOieg0fGQYOtSamfKVprf42sb9FVOQHrHP8DOlBm9DBElgqbmYAwRoBDC62cV
NH/37G6ahn1kxpu9y/DhRhMEM85H5grBFr+9aaVRgxknvQmCeChl+7vkVmMhwBrR
j9rhBSl2wPC2Y2VvqBEDJtAg7EmE2k171pYX+32YITK62LySfhpxj6ErKN/i4bM7
L2R+D3YQBFccqkgtZLMAikjVWszBSmgtHBC99qF/or7T99iNtj4GPJNbRvRJ9Jqy
rVC33KMxz3PwP31qKBIC8auFCZDCuE2s6XbCOTlSN+GggsYczvqxPGFxR9CzM3PK
rWHFsHONCQ6uHPfoAJeGAjQy1ZzFUKKJzRHevCmNTdDeYxfDabSSGXOqJzYzJw72
0J6vdX6Mr9Pm21l86BmF2UGceA/k+vmmPfWSqZtN7DClEjlyKqWNeegGx4bADPlq
UxRUB6w892iUzDzCtsMiBRC9mPiAF5dAGV5oSXBFm9Q4hrEcqLmY50di/aodvgO9
/Rg6Y9a8IrtxOFIzI/d2WL27DGw/RmmWq8+Facgw6OjpLtqYwh7wqm44xcTn+Wo3
BodPNXEi8nuyZQxXpiRkPjG0QgnDUP3WvOFwUJ5c8Zwi1rU5m6ImPQTzCgcXJYR9
OJcOBqjVp5H/Vvcr/UuxPgur4slnlkxSpcAtM0THtsx7X1AXwK/1pn7fs3R4jKFE
OeXAx3W3l2uVX5GGOucabP8GS3N5gsSZ9ZFtnp71Bu3ObxC1HptajhmWlOHZUxfX
z15fS5bT9gYXmyTR6a0Rij5zumItiLXL1aB7MsmTXtkFREU0tzx9EMZFxhmf8l+/
7NJPbF6tKfcK6ajQ2CZFRTlwRxS+h/zVVr9oYMfBEaY2yK1dEyXlHRwik6dFj8cj
e2amWRz8hgTChjFPXPisoTCC3C3MhJxUYcCwofgDCxJfOnesS7PWOgw+JbUf0HWt
BQJdldoKVuBopFYFWhutrV87H4Wg+QHCj59zjDajbG3AJvPocoWai8ZPfJni4m/V
qwOj64PW/KqOm9Tyk+6ijCr0+WjfS8zcDd/350xf1yLA408M0zviy1xrhD5pyZGN
qezpVKHfedmEgeUH6ujxuegdrZnKOpyg/1XU4BUZ8cdQRxCfHp/QUyejAP0jmnf4
Yk9EcU2klnG7MKatdFdYpG1RkxOTu+yQX0prQxFR22Bg41+xZv6ZwPjmaSTkKe33
3mZCUVtVkmX33MmgqQkNSzow66fXcq04fBlcf2XeAQAROE/8/y9225fFHCRNrT73
xqXhGfRqQs0GAYKXB0xZSn3ivwBrsQZRPFF3dUpu5tC5/bPFCFbFOecD44ZKr/Ys
k66vb7bdHJESoq5rFOMLw4FDdWZcXC2a45vVSTKHJE3rfObveCxCU4/BTpQyEQ3G
RP3RNKtZCvF8dIcDsvP84emkLc0RAKnvQCAjJKWRYEGFjimCSkmoT2pdGI+sjQUV
mf0GNbg6O+25qGrCaaRKO2gCIJo/ddqiNIISyZ7W/xFroH9ur29WLrddRuCv4NuI
vkjGK5kYnsAjaMVmi9TPz947ar5FEdUkWaeOfDWuFOBd+Zf882usapap4CdaXGTS
RME6l8E4y1IttWfY+Inu4X5XFwUxdfZxDfrgMJO8XQw12ianWKlmGLZXbyCXsKIK
bx+dG0C9NEaQF1IbjAM3saL0/Z1FY2bBztFjR92KxlGuEZcDdXP50iIwjSSoYxgL
geRNmdFV+beN2fH8Y/A8fe0Hm+qKbNDhiEiK5h8ibc7EqscChfCt77ddwpq73rbc
nuYM3LB3h2M/1Ggn+wW2nlCpTkql8XX4NqfMsWudbACPjNdJXLOal3Ja1sJbVr3g
zXd0BKHM+eYzYk6CAWaGODYvS0PgyX3UqxXCzAmebQTuuSAN/IJ+9MgIEHKxI4mH
13Lmv4OtD9AmjlZ0n84ObADKGuMaTMZjp/z02algOSOG7MdyccY0ke4n9CeRhCsg
dFYw8ZS7dwVGMg8uJLhaylyQxRz1LWMbJ+jfxodAH4AYlqgrg04m/9bO2MGf/3ei
KpJDc14IKINRR8oufVG063FnT/GP8z+pIWav2f2kKrLbormegWzGAOG6RsVSj0oM
OQIPz0jFzDcJGJi+hEzwoAQnKMUTFH0WiGC1IpYPatk5rYUDkoplVtRXDS7QfJxJ
RE+Tge6etrCUXh3uWJkWl0duBuTfQToUvKJlqzCbCvAprSqRLrNhobQW3xiHB7vV
54esGS35VztgvKKZ/PKCPARpJL/h0z00t6iN5eN6qYxwSV8931WOwitvKGOiLgH1
yCVhqktuyiNvszG/LPZTrsv05DWthS0d1S5hkU0g6X5eabTpG9dSWWjSoyZgR1iK
Tbih/a/vGCv1z2imUfQfG/8Xx/Cq+sNszE60MibJLvo=
//pragma protect end_data_block
//pragma protect digest_block
gs5fpqaTLSCxKUJlDiNnjxXNBPE=
//pragma protect end_digest_block
//pragma protect end_protected
