//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
lehtj3wpxoU/Wb3S2DI5zqhsEy3iPU2jF/cIbAlj/zbFlgLUjHfE3gTMPghvH5Ds
ASLU3ASiA/E7r1ysv8NXaya8JxlbThOEnvtL2g+WCcPODcI9PA/ier2gxgud6aNj
inxkLZPIqNPfn9shVPT/NdDRdydkzaPvCSvCab4aqgfTz3WhjPFIyQ==
//pragma protect end_key_block
//pragma protect digest_block
vOvDD3h45xtXLWfkiIdtBwoocsE=
//pragma protect end_digest_block
//pragma protect data_block
zq7vYbul0sJLXLM2GgI9gunoL+tlzTKcd9X6d16pUkMGxRZX9QxauOLZf6nhiLbj
6kJWuJbre73x84oXXdPC2b3N0U0j83pdPiazsB3LAF0nVvFs0RLdH6F+8fwJeCu3
wXfotlcBauOCfagno94y10v45QpAUwl9NfK5Ik4C9gwk/N3gFQl9okKm0rRoEXJ7
3GxBexRe1Nv4EInRoDGdmZUz9DYi44MptGHXJCypSnzjt494jh+Tv0ly5I3Z9RzQ
bsgkxTZeTn6MXW/tTP/TL/GQxiHKMO5E8bZHm1E9FezrND8hOFGSKHb/nAZ4UheJ
rc7naxf3HX2z3nrWyCMQgndcC5zby21QkWXG/w6Sk7EpdWwajys/pZtR5h/XuVPH
Ch7t+Y0FRyamz5aJWJoO3RqyWfFAn9cBWiRiAAtt2PKavRRAz26276T3+ctr7eiD
+4F8crrjwpaYYGnt7bRmtNQbFcV99fsqm01+0Jbx4rYotQSeO/quNUTNoQhYwfSO
Fgn2bQzwcBtmw33yge8V+P153MVj+aZU5MCvG1RziFaOmao6P+hIqRZTnyuo1Fua
U9xpRPnS/1XPlROG1Tp9BBaocaPl2IJX2jfAzfeX6gxX0aPIpyNwDqli/yue08dA
xKNRIDIvzIk+BxvcE2vj0SDugS08OlIZxNojbSTrp21qhkTINQ1NvRMqieVQs+0p
8DXWlU7nu+kgCPSuYQNarzN75/xZJPSOJdYt2yOREJ/v2uwLyTCMu1FoMjkEyJI5
FN53Kyry9qG7gbQWGHkArQrKYAwkxNX5k44Y6IvwrjaByGPLo07Mmu8qLXwh2WPC
0ydtXLHNwCwR9bRaXb5rRU7CGMj18A1UbG9yas4+I7LFCYMwc6vx0mNXau1TqJHF
4OMeRCmQUrgTsHaJvUl+5XGcDkegrsRib/iFCQPXunxrRxQ2P+EY2jw3chQ+MeqS
eQlAxMjKHaxR+tlGVyyqgJBWDs9Zi+YEAofvdijVGQILJmNciiUYvjP3xuKCw2lX
YDW29DpmM/tVXPAByjHH5TNeWhmM4ZhP3ZK3oFOhsfAzuJ93waFtFfLL+3CGsoC3
l0UHjO6JQ9Y0gjtePR/ek35F24ic4n11ldWzrL77WxOL32VD2sOtTPeEuKmpzExU
wDzi3FX828MSKw8qLmV+draZJcwpn9WG1o+aZkugknv2/2l3BM/q4QR/B7F8cgHp
CwZek4ozFYExvIJJhdUEjmilkJWxON/cobSruWmPak4vYx2O6gIQ2Tdzajj2xCoR
ZVfjPjTS/w5L1iqzThm4ev0ucDBqAWscTVRDruzrBELnxejfoOGuqCIxNqSJ+xJZ
XCLInenjgNE03B0lQeFtJ5fZy1p66pRDgbmY27o7Z56jCcbt0HhK5tZTsUqdF9S9
PS/Zjh/2halsKAFkHKmKsIXPCKfZGCGXXKAH8XQ1Kk4MTDWf600ONaDctDtawfOI
t6BEXPg9cmIIsD8PpjkD0ahNSjK/zu3W2kD6FtFN8j7Y/3CVBnFnReooPsMFMnZy
ZEMbU8e4zlLgpeMw29LS2KGqz3yldkD7DytCWIw02A1phDLEZBzKeUGTUCGx0guK
HUoM6fOYENnTR5BYWpBDTwcudXdvHmtQO0MUMeyvoOgp3DB0UYU+lV03oOkm8DEZ
CuhN58H1eYs1wtTPRSrv+0Xr+77zCqdPp3K/4sgMgtsi+WQZhbxr16HIJbgUpoDG
5UBshBVZIy2KgXfDQX41HVTjtpg+LcOIjCNmhS/Rx17ILbcsabEwAf1YPHyEmFqM
bKjfQpn0TifEdupmW79+msxfbdrH5FWgRYVy7IGmwjpXorwxGVaJtXdpXWnNoGys
2VHujhUQJcfAg4Uexj+OLAjcNqPdQlkrl2v0k9oqt6rjUrBcLPOVDjSH7EOYodQ8
N7gpYn1/x8i14p3vvqo50DjGy6eHjIobwLdqEOcVVDTuHWWXKOAiRfuUMMLiq/GU
J3cshJhNrFr/BunyOJHd0QFFBJUyn1aUMUSOOlFUMIm5OWUD6FFzG5u2iyderiWS
HdV5lyKkW6mdMPoBcPnJsWAIxIG46h/z9uS4MrPmhs9o8dX+4dHd6LouQLk4xF9w
CZMlN/b6UCwfndCPDXNVSEng8j0SCZLNXDt4EwcKqQLMpRyLqgH7ks/eUC/YkinS
pLC8ESLdjeU31qM10+P4S5MASRJCHOEQJYo3yl/md//+DXU6PrCBEhgKWG4mnEZV
ZM93Id5xFVAbyQtzCLmSNPj17Aa9dPofsmXlC7vor5iGOoQxxHNy4Kun4mi8w+1H
+P3bylLm0AaDW4SKWz19TWa5344g3F0f2EWmtmC7dgYJZwgu7nvrYs6YZO2mgf7v
gjWErX/TqFa8T/XmMtNukRqXL3iF4rmGb+2wbjgfY2TOO0GQrNF5sIyjIe3/rUyx
C8pMTgxW0ZjkKhmFCtpOZ18zhxRaJDvMUSIqW3Opa3/cfBDzgMH9Y7KdMHS0/4ZP
DdtDarI5oVrc7joSuW2TuamY+8nLYReLflCVbvt70kNlJKLD6Am06ZTzc67/4+gp
YX+dUs+LMQHicDJkyX1C2PQI5LWS1bc0Slh6KnCLXL5ARSKP9IlMnQAsoW36SsK8
aY79GtIyVPzAuR9MA5QWfOdYwYuIPnnQcXXcV0VQWJEnsV4gRmR27cFbV3dWsC5l
a3TR+qN8tSHjbG+q/5ouTNHKEANIVVGUhfbhLP7kOTjed3DIrzgVQ/5DBl6R/BEE
ZPKSYJfpWDL5Vw19bs3uoy8EynFSDfVcGIV3t39ZcoVVHsf3l6rTm7b9sJXZSPpQ
m51Hzo+LJJCwLjulMxHVCIj0WGymUrarp6qZ29e8yuAWLT9dozvMMmMnFbIK6A12
H/7y6uRITpk5tKl1PQnI5xNI+nJ3r8yksRomGnVXqpG/a++5LFf33UIrwWJd5CoF
hHC7IFgSgNoEElb+HVdHEyB/fDm0Fx/MRhV3wuVdTKJqiENt41L8x0g7bhIz/LFl
Ny80x5THPT+dFPu0TZHMDUv4BW23sGjpaCWr7Zil52o4xoEkp5PhiXPNYw9A+6tE
NQYXP7GWagI+nfY5XDR6rrFxIvvbff6WFDqhI3a5QRpqjfBnYaESmEgOZST3pw1t
dhUDJAZlm+NfDunORo89oGWOFNP5yAfGKENwp8SEzzxVhoRBInbmqyExPJHN4k18
gCt2GUaKlU53DmQ83J0n6x345kbH0nCFhZmv4z3oP7GBOJdDmBlMNI+qMrEQpK7p
IleP5OEDXcBA98LdbugkbpKDatdTD2w14qTZoWRbaS2feK2/Nq/TybQLb5wnbIWF
YjDaEf/C6q42g6Sinxtk3SP9xfFszsQub4XoI2S9y2WaQF2YUpqRUN0jl33sjxp/
Bphq/7+EHYNte4Vvlnpy0WT99xUN8aBNvJ04B+byveFIgNCX6l4oPFXCp69d5mfi
5Q6smTpXPhOl/sSag6n2V1xH4M7OQKjJMRHQOgeMHFCmwdR3HyrYfLdDRt/nPUw0
kw1suu3elW3ZZ6kUWg6tvFfUdI5lzYpXwnjdKbfPtvU07VRDNyP8p+SsWYHgcox9
NvxiY43+mjoJrohwQ2loJOMOB41TzrA9dr8fFTU9baIUs9CpKdXu6kqfDIGHUqIH
XzykYMgRho+XoyzwVDwGreG82i/Tpgv8Bj6EsCoKxpaBkPYRjfFSqFz2OamPqBE7
KaC9G3fP2Bq8c3T702ZlIXAwLSdtKiCMQyCAkyG4YBi6TKU/+LlsxahaOFJO2MxM
zopw27aN33j0eKNVlBODC12MNnydlm2jrq3VQw2sF0GsChM7JEJQk8Hsbct/laR6
DDGZQeEgNS2WxBDfDFEcyjlPCHbBN70tTlMHhaYl8bFeT/mdEv1puv99OmtH/SO9
r4vtpUSuVvcUZZRB0p88E0jaXGzICsiHQ0Po7esK18eqe0OMmjXUVfUZY8AKhAJz
qLmyKle3bVgupSaoKp1yzePW1PpssHiXOR+OCdf8IvfxVTzLXDji06ao2aSRy3kC
OuSqP1+MUHz/SHbjxPy5/PDH9pUxL7Rs27V2WgU1yogHoXq4WkGFtppdgBjSmLuR
mPB8fBcXLQoBrTUFjbNG1fvVJSfA3+yTE3jkaGTPoDi5s0RYW3wp4yNib3IxO+Y7
o5bGC3DJuUywiK4xLUwYKHsbH/fwuL8ziIqjw9LYn8d5vKD19RvXT9rM9kAUaqlM
cyH3sB9qUhtKpWiGPN4Wc32jaByUq2m9XUHGD0X6XZX3nG4qGHP9YQW6BnhH7MyN
5VzrvVx6U+qtfvHTXd/0NAgublGs8Lc+KQVlJAFJLQl85cGQVSnL0dffk/uSaNhb
5L5lz3ktHdijy5t4FHVTydIfUK7x98NPFtAJ03MCf1DphUVhP51/6h0wBHwwMD0O
M3XHZnRsak0LKGgRkP54PG7KRCCYYBZBPeULWQLI8oziI9MoB9qzpKViRfLuozcW
z4e1l+3NucpLH47OUv22Mj+8RY1ikM4763xqvLVG0bQDlEMjk+vrRRg4HCdAayyc
P9THtCcFDRoScxHzc3We3k5FiBbRDBStaFmNuX9paDRwCFrLwHxVVReJ6sd6aXsw
yiUjl6A+Lj+Vg44PtoX283ho/F8w+HFaTMZKRMHdnfSqdfOotHYTpXzx/rlvzHR6
7lN0O/vuYPC1HSpTVakJS211S58FTNLBUk5hXY83s4XWLJGVQ0RzhpWzadYJfWoK
exkxOW4BV5+FPXXB8K7hyeizFCVB3DsampmRlkwiukYvwSe590rnmE3se6dEC14a
kYUdtNHM0aYcAkdScIDUCV+LZG8Vali3JqfwQ5yE35fzctQCuWx3Q1j2wM1NkRJf
Oev4bpKO81OxbbsWBBd6lgY7SvnwqKspik0QF/Jqo2Mgiv4y+C786LDHIAAFwPH6
uJa4kAiUbBsqX5C7nGRqrNGDzSsaExRqCl9k6ul3eVyMdMCvuj+S3+OJc+cs+EMF
2DosDnSYNBEdZ9saOar/rG1VE0scxmpoByD2dGnN/X9vrYc1cdzEnFs7YyL8e8eq
KlsGhR39iYMEpqGRjXE1A3gx/EdeNNG1mBUEaYOstLb7wvIKleSBYet/YdReK1vn
5cHkrd8J9fGqzHFFIeGSe4HF5PLAd1fhBn7N7WbuwsGr4I7/uhXVQ05it4UjyUGU
Su3lYrj+XAPp3ja6wprRbKegXSXuK4ANuVs5TLVMi8s7sHQB9x/LiwK7sqeau5i3
oFIUBMqyFgbM6qeIK18E7oz7pv3X0W8PSPJJeihg+TnjkY/beOIajH8B8UDVX1Ng
nb+cRQqMCSi0rxdVdYsEP5osh41UuCDVXXR+1a4l/42KUijZel5+4C3kY9YPrDNp
mWq8vedSUFZZgch1CL7LaEed0iYqs9Qq0Fwd3LIhwJ1m47bn/bHGMOg98AU8jlHp
X4N346dw+/Lf9Mv81BBFejOnUuAT4Nkp0Z1iUD3X9UH5G5Osf0e20xOU2w0qV6tz
NcQcwp/qvt48dtdddGgmNk2lIUF580SOXEmPM06vtkIpH14GnkOAJ7RPZ4pLnI57
ukpev9VToLq1Myn+eBFnYNdEuYpakBFFSlizM25hf/GXii1FKvi259+etkZfnA62
i4y1um0WWfi62SvvfxwonM5Dj2V/Zp5vUthCN9yxe1Qpk8IG83k3XRY2ugG0LkdN
NJL/gz4nB9cFHoSH79+bAA7RwEib6V6RcgqCTB28pv4PbEKShjwJtMNE0Sy8xSgZ
KqSz1uQZZKsrYEuSYNDkvWQ7PqvHtmCjr7HDKSRm2nFqF4E2MTohwWNcFuAokemD
2dR+0y3Khv+IdxpqQ8ITp/Var0Ubm7i+oKIz/AEfwwZ76r1kEUKztLA2K5zz+u7G
y/ChHXJdCMPBhZCj17NG0AXihnVYdwLGMz4TBLmnimMVl8dRNbvz+M8CcdTxc7kY
61YWmmNfVLhVi94RUl8a6nBT3ndVGf+eGPTSgmTYZImNLaZ9I3WmRl5kdl8k1hPf
9myzInMHA6r0lhNc1Povk6/08cmPI+MztumzGrJB9q8C0RAkeYPzlSwXZ8IrGYQ8
YOl3CQzRh4ZPcQ5RvZg9/pJLZyXMlBXo45+dpf0idD1X+9aN4WV+U3kMRm7DWag4
HnnJ7DiJlrUfEbQmQavLMZY6RfSzmn+XL8+FUjWrrtaEUOLcOmbOBvKTxqvjkoXn
HMohMD6XWgZ9ounWiTqM7PsG0+XVIurDUbBiVzftgP51svczFTxFfzW9h2fNTEmh
7tHXkLCri5JVqO2Jb0WkHm2sDFNpVJi77AbALO3SgretOJeqt4DBtPABOdlclb+p
wSO2dEgnVe5BPJt4Vdy6gAZgDg8ZWMYgt1CDSmy3nGA80AiZyw3igD+fCxhsZeey
tq1c7c0oyzKgRZn8owUJ03dtN858dnB3O7Z3KoyOhQ9dhTKtofGhXHcpWYOwiDje
YMfvJ4KLqP7T04zHL0l4cLM8ti/1t/SbmUJJQE9aGrj7l/8uxSKFDk6i0DkOrvUK
NfuGJznFKCM7R1NSCguhl1bjgcNsDl7qLcUpeC6TrYMYJfFh7mmu0N0vSx5ng6JM
D6UEbIrMiuivvqlUQMf4j/HpXAOZ5nVVE9zSlbfwf2c3PL6gDN8AZ2eI0O/I10RZ
90i459Bc6CHcmYdFb0BeDPMwLXyhEyrMBSYHRmHY9NLv6a59pa/6uT84eVtmMMUm
WAH78qbPH1X1Gd1LSWkmag9DJ3ztTfr0C4hzdJUSvTT6KaPCQmCF2aFI1GfQME0I
K6oMRUqAYur6lvbewFM77fmBFBvjHzCu9Jv/unDLcu3WPKEtx2G3JYtv9bo7k8Wn
1D2qTSVs2qg/1Wu00CSzEAvJMvTjYVt9AeimzXrZ6hi5IpKUO1DsVYBTQ8EIpHhO
Lzxpkf+hAe/vne77+WO6rwrgsweYdFsaU962nA/tINxXNd2A09VSSOnYsjNtvHai
vDMpVJedM+VCUnMJxnxbtYiC2YRltkc3yxUCIn45KeXNteTDjA2wrorFvp32zMUP
C+X2SfZnfD9ocJJSdvgB0wITSi4w8ZoB8oAQuigGaA+/34t9/ZtzwSjugnlsYI0Q
4wplz2zycG8p+IgPfhr0d7DqIQEqNXjO4YKv69SzpLTxkT5RRoCfz0ubCarcw2fC
28OVkAjjWkV5wiIAKQ4QTD78pcA24/GOX9F7zFClS/Y4Gxq0TbAyE/ulqeuFqght
fkhXMe1zELZY4oPHX29AJuvxOMqhL+N6Ea7ofFPL9PM07wpebT6h8r3UzYqwdBty
l24B1vAIGbxACKbcjdSgUoPuGDKrY0U/HqA54nT3/+SH51jfiJAHwf5GpfkvNLHc
HH9fjh/o/C9AZC2JTyWJs4GS8PETFktFxNsTldfrCoQe+S4336FkLf+uyrmmZFA/
0UlCHfElqOD5n/8rxTRvUSmIcteM+mNM0pB8smS0Jay9l+XmczCbUtNEezwUIsW5
1A479Y31ON/QSroKIYUEc3CA1xMlOPTQY7KYb8MF5+Kpph/P6PCZ+dWgI2bLP11l
ajAaHJ7WEPznSxoRtferppbu7H/rUJpmUf4CTF5R2HtWCCLcbOMYWi9tczvHEcNF
GbVAcq6Q/b8oviLHjC3y2d6y5c/S8oarPZgV9KQKhYMARf1xi5kRHUI5svxEW0Ik
AWWcRaywGLOOu6YZfRiUJfzZHwcm/cwFtwmSkKFkVoou+zNl4NKwHx75alxBUH5T
hKfsa+moxkYnFKUKLX6F7o0zJRIIOFAaL7TZM0G2BeGbz63mEcswW6LGtV8TUncQ
XT5InNu7DyKmQI46+w5LqCXBunDcpssh7G3R9F0QuuC8R0vrhTsv4uqit6kzgxX8
Nnahv/Xd3J1M9OMQFrbsfNkptyERsWpe6cIKHWR8h89D8eNjJijElavefuH6RTeS
tqK8b/Eo7pySmgJW2RasgLXZEjFsT2uwQI4rJptl5M6ulgmqnlPnmKoaRIpBQC5Q
Rp1ujqYQrpO8fKfiFcExtK6AuIQNPPwpGTPOR+Aih66Pwz35f33+WHOFkt/xXxXV
MR1JS04dygztUa9By5itdTAm0DqJdc+5YmsNq7AbhKL2+ug0wneUvFAcZoB0WbCC
EB6MXMncKOpCXuBVFfJwLhEcJ3x4olpHmYIobyWj6aqIe1JAdsE3eQT1Nlpo9Pqj
k1JKrqwHvXPikFwEtX+YUahWFCqhPopPBG5oHn/+Vu7SM/98RiK/DKuZngg1q2n+
91GSAEb/G5qkM9ckTJSz+h8cVpu4Kv7cKEMi8PYMyz4N+iEHrTGg/MyLeMakWzzn
GNjOaLn77lzuY6zpnZ6AMnO48XkV0AJc/6XYdPBhZ5PZza4kZcLp4U06hnsgCkO5
sVzRpg/zVFk6H1HyWdByKggqhactnyvLicQ987EALEX8KTQ+GZkEIxvqYeiaB59r
98LpnWyEAsWmKHI7IKUDd8aKhAiGHmWzB9v8fLna2W64XNTl80Y2BlEkLexIE+3I
/KhJ2ocdRjf7ozsiv9ORZ5aeKjJneKz9ywXM4Gha6Pi6m7+P9vPlCqqJb64nJy8k
pQcH9acGXLMG/vRUiQ//kqoBgVkmyYfQNP4qJBITsLWixgm5qFxbXGcMFB5q0Eea
LtsgLru0gUhT9RXEsiQ5zWn5LBhhvIKmuHpLEb3VFLg5g/HOgvV7guVLpTkpHEPg
M06pE1K1VjyKAPxFJunDHrHAP76QwygCprmjtvS7YHOf8ZGjet8EGJhGiJu5noC8
RJu9Si3nDIEmO6mqAB9wSoVjIDpuPzvHo+g8eQO0fWmw902Fr9ncAfJPBRjGTK7t
UguwKr9h3e5Z6DiSYIK323t+ghLriyGIYT/BSdLcKw4Mb5BwMeACSr0a/gEiCtqA
5Nji1V1tz5p+3O/utuQoh/604+r9EdJvsh42LdGEK75kdzA82/KA+DRZ0raLJ3EP
630lFxg+KaT9yeaoBR55i0cJZ7VAfKiZ482EEsktrobWr0k0wyCgLodbSeapgEke
osBOXcS62t110al6Aipocbqy4rOgus445xywsBfqfwppCPGlOM14FijhBAxPibXZ
WhJXG3LQbYjwq1MJzO6/a2Bayv9E5PbPX/hospPv4vxp5m3cJ8aALMtlouHon6l3
hcxJzAryqDu1wlvlqvPY7+iFbjo0DxBN2IyVpAbWwkiJoRKedDqZbw1jrLqcQ8y7
Tm1mjewheqlB+Q5DzcGcobYMjaFekqtl3h4P+FXJeevfulqSMmUcfu62dkfQkEEg
Zdod/iXmmNU4nKhAroZtYVdet7BkMBQMUoQZD8FM35ipUCEvMO0d4QsfiA211fwP
fjTuGP5dg0CagH7FJlX0BKZQTIBItXGo07qZi+xJZGG4Cn1RBj9CkyMnTlPrJzMQ
2c6zmS7nMEzgMI512yjgSY4Qqnj9vVOHuRl4Cz2+rQZz73f0GIIVCDHpO3+giCtS
J9l3Uefs4LqdtSkZ8Z3WVqaR9VKFhr6AYbNH2XObA/esscZrWy5NRK0XQXO9KIy6
0HdvgPDJYtCM7Yf53idxx0Yjq4mQDU+UlFJNbmvPyAf6h+UrHns254ILJmv5uxJ/
A95EhJwkwZCqehYQ2RDsIpK8JespYfrsdOxi97AjP48HGXjXa7uIPwnkVBI/MONI
aaLeDYSEQA81XzwwTCU6ZQzeyCRljmeu6sFm/nFKZ32YeNfrq7pyVUvMVA4Pru6f
b1U70ffTnYr0OXIIppBSJcCBHbUd4VxXKzHQlnASv8por0N8jihTXkJ1uIZ2xrZf
hyL+PX1pFZSBb/D1fcKHyRFFU9ldx9GBfVugbQCtofnUogw3y5zsXp+2psovVUiL
2gsjJpBDFljOuxz6QAT4tElz0XPY2jgIc50MDtOB92+HmRLlOCHTwTmjwhzfGwwk
pXCALroQ3HRWObabkXrOXGQDBdXYS2uchRhde+uqHHL+7Y4U1aHCjEJly0ytydkZ
MUEiTiZBo2iPXajadJ82+W5LCUKtHwTvBMT2dsKHTnUIPAhV1S+NC17KeqZ155Zn
GtIV3yIBdob6kzwGShkeZegSIflICEAa2YNV3QFxSHFZ4T1UqBPjrpW6VY1FZyOe
p6GVRjdz/MhIrT0rVUzE54XDZou/sG9HmBemDk8mUkm6L9pSFhX0X+NMrzOiCLm7
aHWCh9dsvECE1vPXY91tJHdvVPSkUV6KDOdUipuEN0qjTCOICHWJyH8EuolmVOKz
z8o0fPmCRgIc6kECQO0iF8cp6oQadaKvbPxjs/Qyhvbdt13PT09Nhd0M+Ut23CDw
oTIsvwLiAn5OhAraMzn4tgbh04IqMfv0Zbmk2TETPTVktutTgqtcVCCV92xwnLIm
XpjnBuCj+OunGsp2NCigu774PpiSoOa0sNmX61PBc6J2/9NB6ctmkpQQsxJlNA9R
6yL4YlpZnEle5oTCnZkkgT54Q5KOfVzmUPNAiQkcB+JDtHxhcNV+690xLTNzUWOa
aDtQzeTn9C5YphB0YipRE6YFce7f+ax0OkHFBsQOp5qjpo006zIpGp1ozOUgoNrQ
NuKSJXt5c4kCwdghGZpdpuiSHYPeFG2mW+5RuQFo2pyu1jj6RR6JgLrLvH/l8dST
IZgikFk07sYSuv4zoie9nohIk2TUVSNTW20VMzc5bh5OcvGft8828p46DPTVq/xH
6oDa4DmEQt0ufoc5HHVk5zk8YsLoRqsGdQxJZspBCIU398lwicFkKR5Epvmx9h9+
izeWD66boqp9K/s8RZxgkBsTawQU6EjTQE2ZcH+KTfGTEbVhOYaZXhusJNAjUEl6
mcpF6GeZb+gS6ano6BmnLpr4aplcAjjl45/Y9z3PPcLuVeLS1rgnerc8dRRpIDQ6
76vAl9iIe1BWqF8j4LdiOwYKNIyE1g7HkH8r41Z9IlbazevbR5Dhx0WvNbKTqaHy
psIa0qj9mFaB5tVorRxBvFHyuNPIAyz5fzE7sxfZ817X+V+7vqt2v2HfQwOlocx0
5hjLJcal6NUEoQIHPzR6YCNX8dAMJplzAupHA23v1jlHBZ6wkohC0TwkEA8I6O6a
J2NYfAafogLpjSbzYc+emuzE1PqJwuqHdt5eilkpHy2FVFewdQNCbpHJNN/Zxw/y
9CJ2AT4n//o/OKfKMu5bR8DFQ/nTZlQDmomqpOOuXMOfWUbMLHLYAGxIKHyTV+Q1
4PyJHRBUz08UVgsd8e+2T889b1SGirg8vN9+lLxnfsvlFnNOTVFtVKYRQFpjpY0C
QTdyqPaBUMyX+8uGvUSOAW0njRQcsWeK3h00NfXqCbBGzjetscsJEO+MWOiY2SGH
1Kz5cC0qYJDvWzhfgJ8CfcaQRXSWTgQo96LYV2sJueWScDMZBEnmQAhOwkoOVyVG
viFk11LPERyFCFDQn63yE8Ej/eF3GC9srrSZOM3s6/+uOkXcVONxsJ072UpLfTZp
6kinFKR+2mrKy5s4fRZVljTvnLbUO6q6+NWU2eAVBOlDg4us4IKc/mQD+pcXEhJ8
s042KRl0fB9G+2R6jXHRgF8YiqTMKMY1mty7Q1KfSPE35Gm3UYn6pKMYCi1y0Sfn
pLv4Dsh9mpcB6S9PDQnVex5GGZO+FgGftSL4bseLP9Wv/zL1IdyusdufgMK/uWyi
fmjYvkaP8EAED2aktQ0mU+0WJV6xxCZJpyeJbuFDBd0wJUIP5lHG1EPJUBb1bKEn
TePvRVbJkgEw9jpD9nGio2UpQ5CyeC+RMU5h5zYJaBfYDvfszTj1aCL14a/Vx1T3
uTRfaaC1BjqRdfBzoSc0TUYRH1UVdJbA4mDfo69uG2Z2zmzjAeyrk9zTSpvLAQ/Q
s/QOLBmwyJ/hiOAT0/EEt9OIGwj+yUkYS1Yc6t6QSOcmv8d13kKCL9tnuDyYZFic
520vvKZfYq5jfx8L3L6xmFao2mRzOTAPUrLvh7d3o6gr2kYRYRhKWK0Ggln+xN9/
mlI8qXhAvGgNCxC4X1wcgBJsTcCUGkqyTgQuy5SpYorBGn38CSB1j2kk8SHkh5wi
q8nmo3Cxit8cVg1RR3xSLOfASaFxL9agjhwiHjhgfuyK76qB2AqVWqdyUq81wVIS
2YRC5Bm48CId7x/qz63Qy2ar+ZQz5OtPhz91g69rAY8AEAXH/vL2yqatp6BR/XT5
4gag9dtbsmHkcED9UwIpwGnhCyPcB7uGJ77d8FHyVIlPQQOY2wBqgYLodMOMNcW8
pVdt0+8oIpfQqSauITFoOn7Pv953rJSif3wp7Ir5rNwmbqPOsEddiTDyxh6JR3h6
BV09GSLKxcZUG0CmyXyw5vhpfYEuyPO8Rr1wxOkpu5GFXWxSHIUJlqp9Y2xfo/xj
vEuQ2eHf7AnDvJtPpNgCSFiN/ZXp3x7Cl1qQxWbFyCU4hXC+p/J5NXIhTDQBAols
/gPAWvxXKkuf61+VGV60NvpJ0dFHm+IwTW+zWj9VF2L8xzI5iWjHeD2c8m3gomra
OkKlImg9LDltKlRbUEc/KuRgC0BJnQSAfbEiSe5vQXB6odM96EtpYfvVbY9/gDBJ
rUjIE7kfPTRxLiOLyq2q6Lt0At0PWkaNq6Eoknk6pqPjpjdpPDXI1ZUs7irSyFzk
oymDSaKDFy3pUkmLhszw5hduv/6B20f7Y4MWVHetkwMtnSfymghg05AyMycDyrXK
WzPQGN5dbhCruLA7rvQUOpn/HuhmsdFf4Sq4PoNBmgQoywac4j+cTNUmoqUQQFwy
GN7/K78jxi/6FOWxHKew60C+eRUpX9tpNpyItgnSeJgU0HnQlOy5NKU6bIsvbcFY
rZYOF4ow65apcJt7j27wez4WEBXBDZ1IeofAHz8cKAyfQuqI9Q2PwucHvZSsd71f
k+nt0cmwzQmTVPJPdMo6cnCuv6MlP0clRwO/vh5ETaQZL03F2sz+6dtMV4FbCD7R
DsccIG8Yr/uK+iF1vBtnEe1QJEIYWsV/PRx1T99BZQoeJQdfIsdCh4j907VkTz+S
TQGQxzorpCtIiZ/zJ5TM0RuqcumTYRql0dcPr/uRT/AHtE8yB54zac9HC5GJvbcf
pSV1WXGd8s+ToasBsVTy8LSB3eWVIf69RtYk8FHIFxxuYCGXKvlMLHhBJ4pk137z
Zq7ojbXrbs2RCJvrVHdaad191ogYNY8rxUORcOJ/205tseIREgffVDS8BikAWQpG
glJllnC9/PVpkjBluysx9hgCeMqX2ec+muLInYNHHWSY5iY+tgNUaXCFEU4HNlh2
HXGgKdGzXoFXQEk29q2FTw0xY/5a+dVYfpY+imbXEEudlzaelbuUD009/8Y9nUvp
w7VOQhK/i42aoewPz9kK0yADfKvyvBiqD8NwaLFynoiPhVEkYoNkMWgQAcX4ZAJT
v9srMuNWqYdwCbxWmGEIVHqokyJaMiXWOrcYh1czOnUsWv3uxECYFehz2+At+9Zr
9+UOgrA9N3xlkqe2lIWCX1/2AKVHHJPG0vKbulQBWV6Ngxcm8+MXIzrG6QFXNQ7Y
6e+2WqSC7DXZhH9b8CbFmy41FQswPWLRLxtf48llM469OyLm3qrTFIY8mxUWFN6m
IiM5mZ0xr4wLeC0OCiA9HgGst+h9K1zlSj4j0RDHHBa7CZjQVIsLj2PeG2p+dnkN
L1EA1JXDG5hl+FlWzyAmDOO6rgN/nv90ur+jbIBTfJlabmnbRdypDaG6pD1P6hmF
0blGZSgngNOoUThNDONAU5VE7QyNFQaW2BlPxAfniH2Y82sZl7spqfkjB5lR8h5W
/8fUEkp6ErFtyH7NxcyPBK33WfP6loNxxjd1+Hot6MzHK13EWHCOMaJxpMmmSrxX
Ah4NAnfsjbhpWHkTiNaCPooHG54bBM7mKGfj8aA7yNHlD+4xIf6/CSltKJrRchid
aC7umWqbr013BYBDZNuRlo32jyk5ixAUy/5UZQjTRxNz0TZAgqbv0GYCkOWBTafZ
tdSfIpNXBQX99RwVXOIkjbjAw0dKAUTQGY8kfWk/JDt3TimoitPpyhyIhC3RzHEm
X+wwALkvSp6rpyHeGdaZ+NVk7FIGcHwPyx1quoLn9pGRBap0rcOIn6qa771R16xw
lP+ctmqovzOcjOfzoGj7ekONPVbr1ceZLTp7ekAFv49yQ/+pq2kCQCDJwbHVNAMY
BERrHJwfdalww+OpCdiLbHu/Q0DjFxtQnuLtM/aT1jrK23jv4/EQNnwdTxmjvTGR
GTTxhTLAeT0yIUCL2g2RVaH9TX568326je5OkZinjaOEUoYrdjBpqYUuZ469oH+J
QRi74m3YjHn7v9AuS9ei4Rf6wozePsDBL+8I2IJl79zdLjKpYaRFl4Gw7/nv6HD/
N2zYGIwvLDNLUnW7D7BjT4Q3H1MWkd6LytLw0RrAIRlG8hxqrCGp0mJ35v3RFGCR
aQD4rjkGPSTWfw1c29xT/bBr9BCnNe1jWNpk8Ya4vQDf+bhU7DQtcFUvLgsi2GQv
U2tMxD6A3QN928pvXlT3wlqj02t3wdAW892Fi8pQnJ4rz89GE6p+ZFhapjgpGKIg
/2KpgQwkrCGj7+Qz5QwOzrBR3AYQ/rLFbsqunmIZBrJ+yai+58L458gadSTrRk1H
YsMty/wO8eICFGm9m1jr+0flPawzAMoqX6BBggDaREqLpoBqWMu1KesoQ3GWnk+g
s27nM0swA/wLjxdCQ2/4GkDGz/VW9Q4NzGdz+4Gaz8LMRuW1/fi7ub3JcLtvNQ1j
e2VdpJCSOI2jdegH+MgW2QrV7x1itdgzhRys81N43+RpBorMIOuHNzNARhQAX8A2
kmM14WRXzoy+dWd0Ls3SDB1ME5ekn+fApyd+zwSZoYFwEfj6UtPu4Hnp6MQ+Ex7h
qUkIgf6mNIIGU8euUXG3H1sDQrDVQrJvjKmbeib6YIvcq4+UVtYFZVgbCGOus3hC
/u+BCyMpHJJ0baa9m5hLEzFTYlrNtv5femh9irPrY9AFYLtigJZF6mKbJdAXgRrF
OHHK0nRKjlGr3CZ4UyAGB8y9cW+11LenQCt001L2kGMQfCh2ypLCvmsAleoAeo51
cIeYIaysZzL0vbbWV8i7/+PNr3hbetdqFPGh5fCNaDyIuE6AtcQKMLjgF/j7sieH
Ww2BLrZeb6eb98oEWLRdi5/+2ou+/IW4qNsihxXB8MPuxfBDWXB5M4Wk4g1D2OMw
XJZz/G/R7Us1Ks1QhSgogYOYnf/S51MehGBSD6+I9S6fQZz542ULSoMejdRo7Pkp
1tf8QeAkT+6kOIUrQFChZEXGKPhis4qEoXM5kqyYiTI5kTsFtyWrxElmNzAjhKt5
53XjH2yCu6hjpcBLS9DLQobyt6Ra7McVy8/G8v74gg3tXsIY6jfmEZ2FTSPju200
KdjN9UygT8KR6FULJ5d+KzbNDMN8jAjVefQW8cDhXzQiV3uYUbLH3xHv7pAduNTO
ePoT9HMKF57TWOkkhyhJ92NbFpz71A9GpIUQNDyE1LwItf9tTobKhLKECP0lJ4td
/DT2dqsFcnZuNdl+RKQdBK+qucUpg+LenA6E4yl8qJKYp7gIVEpxLAH85daawQhM
x9i6vamA2kyWdkXVih9k2yH3bjrJcr5y6E7f+my55WSoy08MVMuoleqLy8tG1pZy
jREUSnT3QefDdGtvHJ+4iC20nW/ifw7b3rrL5oxk4bPbJB3mxRboGzTOm1BFJgX7
Z0UeMLqx2g3gC01tvv9ApjDpOUxOzc6IfYRkFAs3FmJwTmV9dG1fqcCPF4Ku5jCX
2PtCYtmUFQ4oDhTbrW1uPtq6wFrBI4HfYC2a+mEMvHMmtdUc8Ec7biH7YMrxvw1P
dCRDvMOiQbBT9AHRzqepXYblQcv9i8BpFoZ65Qw9+bQzl1RNaD+2SpymJx0h68KA
pFFWnE4hMpzUIaDJXdHPjqqX4L8gXebMVCFSNO8uGMjNUwtzWkplWql0flVnoW1N
qjtXt2zR33szwL+3r/+UvL4Utm3xfzibAu/KVeWN3GaG3mdKBSRRyt10ZISmLlkF
A5vOn0Um66V9oMk2EPjtiGtgeQbrPGtKX3thL2FrX3DEA7DVN7hGuMGSa0Caaioz
2/VffqAT8KnygJ/SEpr8qZSbKOOb8J4Nbg4Ak4hNvT6Bpf3RBztlE+ZRY+QaWjuh
7GuNTqWqjrvDEwDyOx0bAMSq9W4o/xEsEESlF1aNpAg8Gasbc46D8yV9pceSujZh
B1G07ryVWzJLPhb5PEJLjJoGzyZ0vFeqR4eEACj4Il2CzglG7RsIIXqMQ8WxD9p1
7q0MbH/Z5I3x7QMBRZbruDZyBihFEcoU/Pbbu1TezwnT7FTArQcw1rEvURrhqyhz
kx9hu4EEDiog22dgGZ1oug0ypztupNXbGyAytiVgfWvkO5PcJfE7oD7wot/eMY5/
xO7rP5sPk14zB3R6d/9PbB5+Hl/fcVnEh2Qb+9gUa9ChkDElgm1BEaCe53FMsFH8
sWXXvl7fBjlwQIFEMrv6yEJgLx+C/XB0qbWQI5doPADuOqukuw3AKCTGvUFtq9OJ
S1pd4ZYAIkjptTMPtrXq5kj54eE/7q7IUaFtTeEWD1y115eoNQnEyul1sJMwoJp2
krMPcW4JiOwgdcW6O/i0M36HzEUgd9a/LdsNZVXd0BqyiWnvOIHHDsHMUqJFv37K
oc5q/o5CSs8AuJZrNbX0ZUvCMwsf5ntB2ruqatKtpZiBXhhpoNC4wr00xnp32Er3
voZoSoLKrzu2HpOBiRFD+RmXL+WvK8agx/bawUCGbAOKZmyvcCJVf8SvyMetMZps
aq6lcoGIzXPG0kSYeMdhRopip4zl+EzDLFfbujSyDpZqkAQSCSEokJHSw0M2QDBl
4fclNr4sqwl+kLM0xIlvcdRKG4px6cAeKFdXQ6oXgpK3LXP44JTQY9r9DzdqyF0E
B2rBtii9Dor1NBzvzgzVof/pNvLoPf8VkvV1455NHa/YK3JKpeUBBx7hpyLq4aCs
cv+WCIhNfpqRrtHS0b6vN0wuob+ktrxVPunuWWKd9CnIRfsNVTeFcz9RSwae8C1r
lMpzI9b9VdcZMXE52mVoruct2O9D7hwh7HlRspZqNsL64xKrX0XWpHBSZXIeHRn6
CWNFOpNnGwCPMFxrIhtPXQ6QgAh6BAO3FqdThIREcoNDSoCPDY017rEg6QFRjl1u
Vcvwo+TQBrXejpgMCJU3WDrwHIeAuriEcBcjKeVN/VBX70OQqsYTtlFZEQENuMCt
/9Bf2iISR0U2BN4X6GdOtDP5j+jqvTainiLIRNDyalKPDqxomXpCoJ3L0yeqXsk9
Kl/bqdFnCcNY0kBwtnUc2qh8c1hkLzaWlPb1ijaTq8g7JRRWM61dqiwMLiDrvyf6
pWKuVrRk1s38UQEdskYQVfyNxeG9bcUHgny10s1dt2+PcRtbfOzmYbccM3MgyWZJ
ZL4Oh1zho26MBIYS3m3LE3zz8nyqNAJGyPkw5SY6MxpYo/eWs4uPolZhetskRRIs
twx59H1Edw3e2LOeWrCUmnn1ONzaLqpmiNurfEj+EucmGwA5Orv30JwkneAPL+PM
NKIe39XSuFbu8vv8Bh+3aZJmFittcwM7UogKubuM/x20pVppAY3FvWZDcYmN65G9
RZcyqfdrC7szSj/01niGOKrlHSLSNX63zQwXEotwcHN0UFzpc9INcU80dH/rQK3C
Tqdrcm4RxGcfrpWlb8JGrQwvR0r6ncAB/r8iVPXHVRrQF0j5E/YgycD5VvbDJ12a
g2I7Zyg8nPDcju4C3X+24vsjPr/F+gagY4iifJ0eZpKCCeQ0T2j+cDFSgb0FWxkW
I9U9xHESLlUV7E7Be8soE4rMcRQJczME1DlfBFeJmkfTOwxEJOv+xKuXIRUDuSEl
ZDzK8NbBuBRLQlHxXGgciTqfu+CJpLJOEX2Kg1qAp2Vx/ZuEvhB0+Wiepear3s8J
NSIz+Hccue077+cFzp+nfNYHVHbbgA+EmeTxYe1xpnrRIPQ/oPsG8DRdoiQKMdAv
h7auUtAAux4Q7+C4r8FuKuh0NekwNStL0FhymyxoUHdSl1mcgSeZN66ctgei0TqO
fW8LGfsuSp4bPootH3R90cy1ZQqm6/4LSxSAr3xtZIbMrwFWMtcMDUraz8ToN7d1
4CH5oDZCaJa/RiU8yCsIheCu6UcWSAjt0PeDZ8KmVq7e5yQLWxEYRlcMpEVe99Dh
WsWWWXK92EhkGWN2WXKdSQqxCuKKZrVvuhnWgG+FMCKaklhTHVlFW7NmyedAEsTw
W2RfTSIydPA3EBhCLArxaLnQo11KQ6NiuBy9t0BVGGS6Ccck1Z/A1L172R2XSdbI
8vS2Vg1vi7jsxq3zNNjLF7wnRxt041AeWe9x/iTGi+17xcyJBesxbNQvuKz8dT9Y
osCFjTW5+WGV5goOjLfRLBpTn+OtJBc7YPTR0c6FDWFykcnFB0pUaIGFw1WX08ib
kUtvTKCFH3njyI4Bm+fkKb6Wh1EPOQ2DNPKG8kKYKwN0IL6XuWlLivUI94p6w17F
CYPk5oyWIbvNa0a2esmz9E+i9hcmkJZ1ZssljvF2HNcs8xLwatuX5JBss18OtOjg
dJTJtRvpQpgQmgUjNfgfd3z3FMltJImZmsvoAnlsYcwrwCrnIrSZjWXEigSUVFSj
oMqLR9mjH8pY5mbKJYn5T8lNHcz3Kbe9nkCoWqEYnGxNFz/nQZsDz5t5yZKWeCZb
yMGKbyezd24IQmeyPU5aL6gpzGcqc3sM4kC27kPNQVwWWIrw01RKXc3U6SkcC2JF
2cRLnyMIpwBppagSJBhx6MF5iPdXxOghKbcfj1O49nMsS5ljD9RV4YsQwAcTxkBw
G1GW55Na0+rA+ithiDhwHjSafm/eEJUDdWa9zHzCnfS1ZMbjZfjj7rVqJ3qAqoGc
zL4+YNXwj/kAE4mgc7uw3pF3QBDBtYNrmHlqS5E/IAfePHWKqOwBDocJBr8fAcoM
FpEWxQzjo2FOXgud3eWewASXQNvG8+pM4u68qeAqOCj9HaNQ5ubXEfEbh3xmbzLk
bg9LLsRKV+pyfZan872asZ5RtfJrxlzVh4TNF7OC2J8U99uEdSWsjx4eBYIkeM+f
068Sv/hd4KsRRbh56MkL1YZ0Kl3kgTEZEsY4KX+++PWmjKzb0hf1VYQrACMMGWuR
qjoD+Exf0Ov0RfgEVOMovpwvAfP3/xG5pvzAr6LLSIdh8fkkumhM/Fys0aQCTdND
GY0YZNELXttWj3E96iWX6J6dZFWUpluWA4b2YJTVdSNlYsjwlIRmJ5x1qr38YWwZ
Wg2g+MnfLy5Ysuh85vi3bIGTbPFP8xJjPEqrIsZcZRHB7TqQ3/F80uKjWSoJyF5i
vhUY7wtBfH5D07i0/Cwz5BGGaUXX8bSJXBuPEILbLH5rn16FYNX0598u7QpPKUXI
KmKsTrBjc6qp56bsUCULIm8DLGB5Gr+DpZT8Ly1SSnToFpNrlkUbHxsjlR2RCFuZ
IODwXaYGx1SRJ0XGjJiNCiJwCJ+ShGDJDjyV6ZqXVN3jDr87tKARGQGrSvN115l0
Yb5MnkXk8fGdPzkKznP7lsou1Z3yJD+hsUmAZNxx63CWO6TmUI289PSXJSbyGF+x
o719MfaASB4GumVUyW61t4PoZlUfxsxKQ6jyczP8To8USx+4PR4Eg16Rapxhe6Yv
pbySzHPWxZCU3AP0URySivHR5yGkgasemYgaWwuniwnLUqMb7pGnBRItd1okS9cM
VRpzqyj+6x9KZZf6rfLM/d35hzJlswJJSs2Ny5G4tJCgNzKbG0nGM1O3yOLH+8cl
31+q+EVVf9IVKSR6M+dzHy7yyiEEdD+rKR7HUgRXpQTibIgYBIFjLd+SUKE9q/a7
d5kyYJJWlkl5/5iR78kfCxu+TpB6ePapBw/QjgQuqHD6D38o6Ox6YGahM+FXU9g2
OL1/86fN0XCr+PuN+62I7HLXAGefYZs4EYJeNSPRujtSZ/988H7FaIxJdvXZgLOw
UcNSdK/SgiySbZ9gG8RxigStg6q3dMAep2QdWbhGeqQ9Yy+HH9ulX/Gxmnn4/Z4z
8JxsAX9SSgZr4au0i9gXR+UxcMA0UUgQLHYOqp7WyDYj9+MJ6mhwITc5pezegq3i
JnvZtSkMJi2ZUATrEcZnQSQlmIpdc3IreVmf9vIEGilGL2wbnLUtXTV4693kqlRQ
kBYvY+C4SqywXn9pcF/SsTAIWZuWaizwEJD5MgEgWbJV9nHe3cth/CUMUn03drp3
0kVBqlOKDQX3+ckPWHtsRNU81IK6LGMONNplCG+fOORwLZbG3d68CV1yM8aqeRSY
jE234loy8l6SEeHrjOizxJjfAAiRPZjnwRtXVw8uFsClip8CFGtoJFdsIR5x0CAk
BAWmUme/4wYACkHTqD1WONlii0oechsVkEZMflc4236IWD9Ceaqv9XjM/fbh0coB
r2vmKXf20vdRrdBckFnIS/7pLEdnJuPt1x7Zb5LpTmuiG6hBTUiyCqTLzLWqQ4Jd
Ch+CVsJ4B33XnUcEisYlLmKtVhY8qOG4HzkJi1MeImhFidnDEK8k7pa452lZqaXu
xkPovWTQqEipF+rVVuwRR1lDjsfsMOyUu3qCHXtA1wQMDYymHHuKosqf7EL6madb
xUoIVLbC3M41XfOkzeJDBUo3P4zkzBIDLeK9IuZoTRN9G6fj0JX7O0u/HhgMwaA8
hFIjKeEw7SvcICtXaV7EX2udra6EV8ylTdwujcDiyPDuhycX4OKAG+o2YB1y37WR
klsoJb7ut/xjxAtie2nKmSxcnYZRu8BQ0xQ1fimgRjygdZIF/xZ6wB8mbwRts7DQ
5BhRCnziyQtdIr9b0eF21ZidjOnjhy0RG6Iwy7Qm/dC8nj0vEHwbrQJHdcdT7avi
jur4RooyOIV8GbeyPRwoQ1gt6esW68Jtc6Ct+DlOpqOcl+IjRPjHV5QGWQAWGXRL
M7cuyGCRECqd6El3k82zEamvYAPSi9F4LA0/0p7OAI5e+McdU/oiv7yileF1zEBv
nmS5A06c9k57ztokgJdBzsajwUYQtL8QBVQ1pBRjYnMJxM8oNvtIXc34hdkrI/6W
9rcNO47YavqdvfSx4HnQ499ds7+xydpH58bZM8CqTgECNgMxLYhFRrihucHZjeIw
aglmuvh4f7HliSzi1yG8Luw7Q+QHqnT81ZrrPPTGfvwsItGunQaYbJlorQEztAoD
32f883PuBwEMWq35bsSQBqPjIh0YEGKQ7+Pl+KmfU4+Mn+ohOpjjihkekeuL2Rqz
LrudYM4zMr2m4c60uM4lHcBm99fxsB2SYVjWtcF0v4qFkNQwYnZmjNcER4Majrrt
FdhJfMhDZ5iWKYJ6aTabkaJ4QsfARDkcqnY7Du6MYxq14tzIRsVQdVwppz+jAWWl
JzUzuOlwPAfL/aCKItfUyPEEEIwmRo7o9TJssVTRWN5FO/Eg/XMJJmOCHBb0jRgO
6eM1D/YnXuUOYxZJxKk+FrpTgESv3h58yaS1Qgz1XgBt6ax8PSfE6n6O+onb6OJs
K+0hFCS4n1GTY5ykKR81bvRM5ZXuzT8m7kktRMKNkXXxj3CpsHc63IGURNFyuHv3
t6/qW2MyXOOWiWtERMaTUK9008ZUZ4szhg7vg5nuXH7MjVTQ2UKBb0u9s3oR8ANt
CejGgBysbLKugp8DxkB5mSC+1ZVJMmG1wftaSMhw4c2+55V3qgKvyHQpAK1MScCu
woj5B6EHVouCMu3fxFp8QPxLO13P3sLXN8AescuZXMxstIURjzoMKxxtuXsTeTlk
rfsACMltoaCpZqYf05PhkXvm3nBtMjgADjZub7axrigpJUpOA9M0F1BNLkewWKMx
oIsf8DX8hxhIh+2rS2dR2yvJj7H0Esi0Oyy5R+dYKHGBFFuXKcs/FtKWrjEEdq7E
O+o8JH3Hidahq80h2UO/ylApxJcpf9frJBEVv5KqCBRZSYu7ncjuxL956EdjBt0c
Vks85uZQwVFAziJEVVD3KS/jgy0HyZy5RILkywPlTdDZYPl4kV+EnoHDK9QxTOFR
dES40W92pKxHWPjrbEp5FImjDCOHXvB1WLrqXZDK/zfxfO//CyTDVhBSXgnraGcy
Bip/6EqnGBPlyMYOwqGjkJRNt7Ncdb6btirJtZ0QhJNcJfwng9cInbFvB1N/PIUQ
VChYZ1U3oo2mrG3KiZUf3o1JSGVl6G95e1mfvL0zV7cYS3mBYLIX4+wclT2Xyla/
JPh61ji0lF6ApxkCpJ2x8pgv9U1wSy9pd0vbS3Fhgld1IM1QraVPs1VYJjFSrxxa
PCLsYaU/UF7HPoPL650GmkxrFj0J7MMqrTEJUVk3pJi/Fya5gdNJd+RPqJmb3tss
Cy4Sd7rVBxDk0bvaQX/FFXFhywytQ45iwjteqWgtWpaSXDtCue8+PRjWjIy5Svq4
49LyKyiVGSFNx0rpxaCuDAUj2aE8MVfmfhU0eNvwcEWWj8dJNoBBtuVV4namXOMn
3Fy7folkggobKT25iBBWweed6nzXxs3SCk68oWMRAew4j61PU0kvyCtBPFFqrmkq
SujZASB+dGXQ4O43ZHlONORXoOYR5rH9pSnwS+Hgngp9YtGB2ZFhiZee+A6Px9dt
krpVweFanCRTNxUecfUcRYe+Izi7l2NcQwp7XLZ0Y0JxxiyJ88oK2lYPl7oYFM1O
uJVKZWK4yEmB7vbU8tJO2GWx9kqe74NAIAg1LQfWLAoVXToaQqN2fQU2eVf6pVDR
seGZTrS+Spi1w2M1BKrDuEGtroy3ljyZ8w/qVT8mZXe2MU9p49TNMQGNnrLjgnsr
UiYoHSesKGhS2BNFsSLfzM4os2fdJS3KKoAuHbE8HBYJCc+So6R/tApDXxNVES0Y
LwYwnkUFH7jOmyTcCGng0icMwylXqx4SdLLZ85mHyT3x23jwHF2Xv/VmcAfpFaYx
mc8vRYoi29pHLnyGJcA+K6ehYsgX9w+51fvzCJAJHCY/XAF5uDit3p1YLdflPt3j
WBDMYjBh/0VfFYbSOd/59H5UjHWPa286mgF0yDilToGDrv63Q6vU4IGurmT1hxLf
Zqh+OwoA8kbrMs7rrGuOg7RJg6+lPnVDwydnANNeVFQpIzjI4u+lD2450YgvAlL4
e4v81GlrmhAgzcJmMVNg5ZUGlVkVUA1b9Fvm3uTdr+tTvp5sHINjxPf4q6JhhP6u
+4dYjCkI0WzHOX74LNV143kF+8PzC8pi6/PrbDm5nGQrSZKp+hRiaE5m3PBuXwct
qjo+aRe1t6Y+pgipbyRcBz/Tuha7RQYOny0qE54z0tSRzDkAnogeDA1MfkauKRwH
YHvF6fiz9xuDcJGVd8EuVG/hnRIHivE19iOJJO80iRJZ99pyu05OZ/nmZpAMFgD+
id6oc4w2JG/PkSthsme2p8Ebu9FYwBiNVdK3KeormpS7oIJP18KCfl9ycbTUVRw1
5anzz3NDymUg+c8yNOuZbiQix/hCo8QthozLttOo0QM0FXILVtL7DKVVFg6mUP36
+y+5XW0NrXmsLqDbHGcPy5LyQP/PKGVnR9IMq9NtOfD8Jz4vgBOrgSPhQP2GgqYH
pahixZzfenJA2bZzQFjFHf+Vdy22DB3jlkI7fZur8baacUems3D2PPBzKIAAkZla
exAXJX9Di0qcT1RHSoVthglylxfsFk6Hzl4d3GgCTovvq3XT1DLgxu2pez4cw/c5
xADywq+YMxmjMWrCOb8z+JG4NfmCEEA3yHaX3Rewf4rEACupzFT22WfZGDq1D4f+
3Oa3rc7t7AwaT9GOEKvCN01ETJz9sCJeh19a1Dn4OzlUnss3yMpkvgkRBUctSWQm
uyddVZA8A7MGx1MyCGYXR1QzA4XQhP0QvzykiIeY2MOlS1Iu6V0XwaXnb2X7Y+zo
x9KIrfIYmkDFft67uYcJeL8ssgrIKZ+puTzUt3nzxTZI10/KStqrWw3RQWSRy7yk
7lQl0OeuInHLMCZZ4U+IJAw5qpFv/oLSeKNuLEfWZ3659iH3VH2X87hCHJwLnWyK
kWP0cmLhZg1VlhWmr6pzsY+HPs8CcXlHgW2/ticZuxWxNx7x1WE4vijISXHOPFbg
rYrYXyIeFnrq+2VsEBGss189kqi2vjhU84OlzTb1N4pq8Oj+xucjRTJXYYgfkAmq
aRN4+S+HlYNXwvhqPU3ORoAqn5Y4vxOjtGxFU8usFe/dQLHtnGZuV6pcBPUsiQMy
nA3G35XHwBkLyhD/Q86X9aZX5BZaZEvW0P37zeJpt4nL8+qeoO6cv/T73RkR1mni
m46yEx1jpB5dSgZK6qjzPzmgSUgdtlDXU5tjHPeSahyE+ngUYcuJQQ+b4wcMYvvt
pEi+cxpJ2yCshtTZbldPyzXCIdujC4CslseZ3k8NsZpExk4AkyrmqlIAK/8uifGI
KgvSru9UepeajODKxk7f6B93+R7JNWm4WlENMqJdzW8FAp1F19mQaX83eqCbyW3C
KeSFbYYYEVTJ1iS4gGuxTny9GJdkcBIhguGJ2U5X5zomHnrfOXY7WNxC664zYyh6
tMHJp4c7QnQaJNGEA/povrzm4IfU2QnTPBNbSm3phIUruh+1+gnn7W9RgaH7aXvk
ZYi2z5aV0tsEDFysl8lv+qldnkYmOWuu7T+77POXJoMGpLe2O90xg26TcfkKEr+w
wXNTH2meKW+jwI+cPgjM1fj1jH0hLUBKNIo0/tHuEFsFeruTK5AFP3fHIfHwINfP
8Kmev07+ojJfdgBJBLFYMXC9sTV1I4Ducceedhfs19mQGYnd0r32i9Bwwye/vt9M
9le21ktLJcxECsWIw7Qn22f1joBsPwi7Sy7WCtlcxjc3e+kYfQA2e30tHST1EARy
jw4eBd4K3WvDmg1thrj07ky4hN69b0OoRZw5UZVAMiuQ+SNHRX8f8YXb8SebM9f2
OfOx6Oof/u4BqXy4blFVlC+7Ob3goL0WCgn8d5GmbN4cSYoBb9Z/3AwU7JWS2dIr
e+PNNRa7eiXLSa2XANDSDg098rswlxw8awXOhGqxoSvwelU5Z+l1B6dQ/yOrGoQX
GV4mmPDeueWOqxT/SNElTgZqg1Cu71VJW3p/92nuARsxb0O/E8D/z1Kh4xGvKNi9
5RUPHJV4LnxojXEjWDXHms1zU9fBhKOO/8NN2RiuRhOuck0dGj4gG4/d3AtXakGl
6V8RnjKMP7uUxlPjk0bDszIwqUtRUXUk4GShG2BsKznD5YdoxaVfNStvFtgztZI6
cFsZGoDXSpN01lVQ+FaYBhnLumHaQE1z6hXMWsSKBtt+wrndDA/NNSr7BJx1zoqD
9FOULts4Pq9b6w5OAegRsBNwbnp7XxELF9Imo1nGcILii0gq9MVp0V4FOGWigyaZ
p3hsDWPciL6MLyqMH3MzBy9ulg4Mi1BzSjP860IgescO9FW6In902iMwEVwW4Eox
sF8IpcOJyYd0IBG+qdQg9STVg4Gg63oShEWw8jwVnEYS31I1VHCd0+RyTaKu1/8q
9t1kERlm15/UUrUxMpyg6CYGHFujPPZM/JnMWLQQ7lKpxaOFXhooMZgFYn6rQYkB
sBqm5SCoQMJntfjH7YyUr19zaU+iz+6kuB2qkF8gs+AuJY1jYFEEsFKIvWi3aDQz
zjMqd4PE65B7LJmZFgW9iDYdi4pZ/euUcMXCMNEnIT+ZfqjjlQk6kNjBUoyKoyn8
A0q8KUQs9ruACLqWzwVODt082Ldp9+ObVdokS2X/f1A/AallQ6lHnNJgnndeRVVr
6E0xJ2QR5j+VOD80/PmnhLKaWhhGuvhexnvv0T3Xfku8kcBSFLPpvkyk8tocYaKE
eBuMiJZ3huazji6jW5xUaDebyIrJvEN7cPALS535iPyNWCs6sLP0EwlKXy5FCWFG
1XIbvi+FQ/o4/AB0lyJGN4ZXa0LEPchV/EK1J9aYRLaIcnhqit7B42qLZ+qRWGaH
z4+nu/vOKu9TSBzhVOleqHELqAwSW+FTZlFhi8Z6aSHPkdOfLwCUpnXzxvW2wdh0
b7l3EGESfJbDRkERHBzF++o6ndkfdCCYrbAUukidUh+pA2mHTmU++IV8qykPIX1e
e7pYPI/JQ9+aJCE91NtwSpCq4/q6hUHJxU9Ft2NYoLY1Wm4E6laShVXnCFD4j7l8
uwkw2Y1JEm5VIR0KVSZ730tDlbznGKVCNjb0nqAA2zytRTjCIloCTzfSt8afMq+/
eUWEzOOmP3qSDByeKEnwTa9cBCVnxy6yD9Kx/fPBqtoLBGFKtH7JvyLPuHeFW7Tu
MqHR219bzsoVYtQ1Fc7UDEpzh4+7+OMG+IaRzw4Bi9aBwO/ytVC80t5jUOitPCbQ
IEhTqDGHwwL3rj9Nchkl/8A9kyXX4hERqyZzieBHK4iLMn3R+Dc61QAhEofmeWis
UR/kF9AEGmS5OEcOVx2fkUbmfzWGGDzoWOvj2JPJmk9RYarMIFyIwA13Pl3pAUPs
aPWHXEzxJYoebKlcHFWqhwiyAtHk2lJht8e4H6XKl0DR82WyC2zEWZSkU4/RLHRC
f7y8EZBA+DEslRlIyCfKxlDZ1TwDkjMliz2rc/lf/S8b8RWXGzCT4z9wsztSihZU
G3WVy77EDYH5xavXBX0xGAncls1/be32JUuJwQhtS9hLx/Tfs8aX59+SAo4Rgsiz
DLljyDGt2pgdqt1jZjW8v+71AWedRSFXqvbRs5UCowv8Rr4XMUlG8RSpBuVhH3et
wslX0vaxo+LdQUZEPU70cKhMBQ0ClONynS92b9TAbBXTzlL1+QIAKhbXGt/WmusT
RCDOEa5MgCoYI7z925RQLfWtYe0D9KJgq06fcG4qlxuNL5XtGGiKAWdHRMOL5cwB
VtxkFdyKGkc5REsoCFiQ0cmRsUI6otmmLKykqVkoQtd6oxlthRYY1x+cWWi5JwtC
nvvioyDiMhFFCLuHfvQKgVUDaKDD7SByIryCeZ2mHa877XkfD0rxeOiSkgiZMjQK
k5LLFq+7Orh0PcC1KeIWWfdXply0wCRizZAK8Zsnz4jsC1lHD4G5FED3d7SULjXf
lZQHc/XqINFRE6zyojkMYTlKt3BRn+dYLMqw1u+6WyaMkhHoCcZcNqWR6P2DKxvG
VPI/uHJrgrYG9faPxoOUTbTIzXJWaCtYwMzj6Ia+tK4EoohYL5GW1vrObI4gN7gL
NmgCnavHb/l1lnVaJ7DfccQS0ShwvYPb+kImL+lBSnX7OjDwkGfKj8ogRZdSUAXZ
Nd5iVmtEdACBPewPh+QPVp818fKNz7ovgbe3r+aTOowCFSlw9F2vW3EP6ZYqGxtx
5gUcQyKM3U8yF/YMBJLCLboUYM1gnmocpRwf05VGWEu61tS7a4GbaddUqmncMxDM
mzIBHqjh/vgwTy6oSDmQbb9g+Wk7mxTTEqMvPprJs+WsjTvLq638VMS1WQtr/yhK
8K6kdeSDXNj6TVyxSxDgIzgmkvmLI7thlZWWZl2xS7Zuhqqy9fUZNIp/Mc1yhCh8
MILOpfCs3M1YrPh+QftiArR6fhhoeZpcfMTrMY0CPpVE8MfYBP34R0Jjcv0DDNhB
oUjHGcUGxMsHvPT4dWvBjIlWOzMSdr1H96NL1Xjm9vWdR47DAMRqD2isM5BM2B6r
1uP19lBczmL1q52fyNL0b/fq2nfgpOIL39BBOaHqSxk6t/ndBy7VAewZkjV6f7V4
6kXowaC8Tu22B6snlKqL0bG6mG+S/Fmu+lkw1nmTGLoRM/Hj+QzYjKr2m/lSNuaM
X84PljpaOfv4y9oSuIEb4IIJwI9YVBAPTEWv+nD1aG+UFpHNaP7Jg75Ey2fYsg/W
RwEA1wTqan+88WTKxMPY48XlJi+A4Jn+ilm/xtx5MbSOGEqSQKGI+5bree/mSW7p
6IN9bkGDbqE3NqUEk+sUt3Xg512psj5crbcJkFYVyLQPDKCNYzYhQ18DgjoyyUHc
4dHEiVYYi8mrSqE4QeZfgTdNPLd+Iyutt7MnueitORDmIDVbUPTV6h8sMETiZviT
CfTjvdKkM8kvYtc5Rt0r+g+WtpoovYa9QrUuPA/ti/+xMI9ilJqsy98GL43py2LV
I/MoQ27mKNh6PI9uHS5DB6+NhJiwVFiQk2f5AJKgidqnFEGDaVP3m/oTgqY4+15J
IV5xEElDsAKnwfdA7P1vQYBZOTXP2SvMj0UF2kEJgAZ/xXs3quOHR1b0qhYDKUFU
R8GltGOwUjK/cmXUYXrixzjy0FT7MRS2ZgBq1V6j9QaR/gslPiVmXyNnU+ba8xpf
IkK4Igh6O91LR22I1RI/Mofzr57QEKAP7rEcKXej3RH1sIMyGiqTGIqPR3XPDQex
vSTa7ev75JVISWtOdSdSYpYCw1ecEwMpob5zyaSJmbZwUPbYWtKBRT7WQ6jDl3Yh
ZIL9pJ0suQslCO2MO0RhR2T4S9f3+WviOmw5+VmGkqCI4eU9gdlZSNCBlUoEY1Pk
O8Z9QZJJPa0u0vgAcZHw/IKxGJ4kmT/Qd+n3NPzfbweQ1FGz/pYH+N8K85WCMERX
ZBc88dcVHUd+kYsQB1mEbk2WOYyho4Kb7dxShOBei49oZ8AVuWzriUzmS/CmESOg
5wqnhiqJtvFT1sEBrlnQwGkIPZmHsvw3apDTVClkLdnYgzfzTyYKhGXefuJoUYvw
l9IJbssOuRIt3Doo0H4abrsOe/cZvi57rQcqYnwcVoXZk1cv/D7C7uzJHZnfwWgJ
GkQFr4j/SXMJZr4vCvhYSkz96ow30mQATRu3D0cAm6DiJx/om+nyr9DgHfAKxuKm
wBzhc08zYXGXnwXykeUu67CzHr1fxJ8Hsoc2dSx1L5PxqzCaJ1lhgFmOKtf9Ouif
K3KDg0ZGimGGc1l5RkeYedoa711ehtqdgYigdbxVCQ7ytdIar4mzGxasIcYYBhRj
eN0gF9J+32fvcUNCY1NaVLlwZpoSdtvb0IxGh3b2MPa6QOBUyNn1jeCLtEfBIFPQ
tESoFteUmztQyQV0+IV7jObhpJwTKZVrGkZsb9EThSDTpO3fTk/4SGhPdP3PnkMc
n4AnxkaVBxB4yagBULlKHKawLQ4XnX1atlqVHs4fAF5NRzvWwzemTftkx3k5emh3
dRprC7hlku7HsaJ5yEXwuszKPC1WoTw4T7MN1rH+fy/zeBJMQvRz5S3kN3kRBrQh
0MDz59nNnu35BCTPAsDhzaM/efBfRQUo8/8327RaMW2C1Prxi/YOeYSUn+Xb+dBT
BGcD+fusWso3x2mSJazVMYb5rk0Oc74G3Z7TpgJKgj+HqMey0JqFV4947yZILsJp
K6QFBNu0KuEVrzu/G3rZHKP1TmmQZaK6zO8GAO4m9Pxn2uIu8igx73LSBJgLQEvH
Q93X+2X+JxWCAHKHhOnOapBevOeO2nHmP5PbW3D7322cjjhqNGpmKz+4+jxlUDhJ
pvKD63lR1TGebnCN50Q3nO/0MYJkbHSd5flTd1Qtk/Usb8Tr4FDg+qKqF825i1n5
h9MIm4QeYlZWWhqecHg6/XsGiveR89p3NhlwLb2keL2sU45mpQTHo1U51JL+7FWg
07/xXGCbOBRgJkuyKKOIHsV6kGeVLwx6cLd6HBDjfQssif2Cq4+HHcx++kv4fxz5
HouMa7o8GYSCgNaxh3lG+aqjEo+GDVJeh0oxMTSuLZfCG82HsUUG1flo5L1NhlZT
6NAgb/8gbr0OktZCKKmP/DcO/YWCbyfGlOQ/TIDOqcWJ9hvLZ5qpC8Ajq1yc8ER2
3SnnQJ0Hqqu+Nn6aGUbFQYTUpGuRMZVLsw43Lm8ufMAVJXFVTTxhx3xeaXfiiXxB
h8EsPsunk9DhyivApDoBXu27y4F0HyWYGWkoirwnpUZyxXioSsWU/1K0GCfHgZit
Xy9ug40r2uYqeCgUApaL2nLryFd7m5QPABhhbGxe58EPYv73inW1TQAqiB+7i/t1
Jbjb8kAhY5H+25kCX9Io4fjkaWLnfyFWnZK8I9dPCiyOUJjPVYuacVmPcW3nNn2I
51JkxWSPZ22sPF7OMBS2d3wAXP7vkXevK1is1qdQbdlN2a99pxU2dKQD4tB30zOl
kbRp5tzeTU8XhfVu41+/2SPDEgDOqYh2G70wcN0W/a6OvdkC1obbiULV5ZVnWxV/
ErpOk0M+5L4aCsBs63XsqVZB7w3h16QT5/lbMli0OU8zVex9YlLi5MPq6JlkIRtj
NtDHa04cCxPsOhnnT6xKrOREOqTd0HALtKjrdD2z05N95Q+AsJ/wcye3pE5JEPID
QizMv0kq79jeYiUyhjQzBZdXb9K+bBLVbTKJxKupPyk+MDA+rql/8NFS3HypIszS
RrtuD6311+56uma46XwzEW+TQo1z/1Xq6br1QdCZ+HT0ac/mV/Z6mhJIrRagE4hl
nkgZ1khFGWMuGcRc0AkPEBaTdnxBh21rHOwdlK4Rw5hRM5E6qQ4/6HoaC7zgdd4j
XwbwoTURQI7tEfexaHFIfL6bWFVvPtlf7Cbf8xRATKYNEECU16r3+Ur5s2hIfGyq
INxZTYrJeh2Frgh9e2En29P6nJjnYMOqa8y4GiJct5z2/rRrJnyL0Z2IlFgp3TA4
0qMQU9zbSTIjTjG9s2V4Y2PbZZt5fTCCYhEI6GrFXcg1nP+dSjCdqpLBgW4I1fCd
xv5e3aXkMuU3tVofxh6WFLxqkpjUYKc6nW3jDfWE9Z9lx/kNzNWrFNidTQCO9oWn
VYt+IZ6aRZoknnpYwqkqMWupSN+ep5R8MYfa/3yR5KBIaI8Cq4tO8NGVGjNimnPE
GYEDeujCKOn0Pk75yAvtDwV0F6h7hGjXpF0Vw+/WEQo4YyHOxyPGUjjCSE8DQLAk
BhaMjOezVZ3IKo7mq9U43oftomg+TBtvRcx1nEq5oJ+x7ZsglWugF6myTPAp4k0Q
EYBZ5I8EUPoNMjURJJ5x3E1HcNRndSEot7dEsC5BtZnEQfzif7HmhTeeJdyqGTue
BKXuYmD7Ytc+W1rJ7sH/hR9OTcWTlZhGQlOJ0keerbbIeGiDwpLpkovzP85L699c
l4zYPI+elI3BOdiM1MnTqCc3PPsf115+XbCsGQPqbIidjl9tws0wI5tTWaR0OS45
jR6RFUAY2wZ9I+q/lGiDl8SUUEbiKnjd4imHYVEK/LVaao/KluYntCxr0tdamOPr
j4oCSsiu/gtJ/XaJP8hD196hcjS0FXQp2iHxi+oPuMlqJnOcqzYEIy5rw8ZR7lP9
RCx4fsCq8Cle0r54ig2vgB2Z7PmU1vKj4K6r/lkiPC9jyVx6E5b233dmmNdWF6oU
aAx6dQ8KJicQJsYxEWJw6ns7oK6GuYygInOl6jxCB1JbITG4azs0IVhGFzbOVwSp
VQBbAORrCzZIs7oQJuMHQcez7e7Ts1K7wOsBcXUFl6Fhuw9WC4PwElsxhppSdfcl
w1sUCWpCn7PGKTidnBxMTU2F1HpLrsfZy7rLTAVm/H4+LDO61kTYikUNxgDFRZ9f
LN50kgw6Bh7VtN+cyxmgyY5Lb2/HWp/U9BKHDxzheM3he0ZI4VDGp4jm+FERtVN5
+TQvHKBNaayFhdQGXOe2sgMenex2NJITNO5ALFAjDHp1GdgvnlhZt6xK3dwLiY5x
3eu4EjzZwiOcHl65deNbZAfxun7LIE1TEEeB1Nk8we9cnHLELnCMlnMDSwNsBHTh
cX1QXIdZQmRTJkaPAkEtRhBlUs4bIXWVHN1htmd01qjDO4gcoB8WkqyYTZ/YTtg5
1Yq0oEkfRzh2XeCNar6sFTrkfLWWsmHZIDVSE12/gnyZhcIvl5P5OSolU+91nG6T
OlSRNcYgYf+9w7hefghsDVY7PlE4D2/6S9ZOT4r/5+/uP3cFkFsuASzxQ2n7Rz2j
VmFo0GS2jQISFZ0CP65bJdCfL1nMaFaqlaWSqSGgm43yk/svUf3Oq7Qh9VbWck8o
36BsKL0Ep+U1A1MkxOR3J9ctTtzZhadFPdAoelyYhBstg1vXtIyNwq7eTH5EjMds
WkbeD78e1WkahT7wSGOxi1wnEgpazXwifgRb9wK+rZEVqDzlOrWFztz57N6By/DM
esyOFJ8shO8LjdJ0YP1X+uTPM7siRkSbrRn+qJosrl0lX9A8AI/+gMXB7o3mcpGv
Hx+q54Fm8dRK0vvBw2ExiegSH2y3cQ7qVZRsoMaIQNgataapSHXRcq2E2vJGeyGX
UaPNCHvPmXivo+Pn5uBYwkw8Fl4ah+lH0Uwv1+lwRdagcm3+RhrZXmfscaxYfGgo
rgtuv7Vd4vQ4p6s+uKvFTbPHpipfJ4A8sRJ98loTglceqBc5IVc9XtgFepLL5PFb
iHNyKfia4z+m4ivxUBXUHK59Ni7oydxCKo+uq63SUXObMQhK3xD5nZq6HD+Bdioe
9uu3PL7xoBElkC3QNvXTHC5+feRyDqv55rTxXsN47p6DHqNNuHBG19xdbTrk8ppj
0juSFkQELji/1FMSKonZotf1bXqblc4NK0LqATbyX3883OW9Zd0wYt6UwrGI0eZS
csNIkw05qHNrBfuMjW8w6nBZwP21pUo87gJ5Nvtwxh5830rQrrUVZpPADc/a9Dts
Q7MdF0IBMh1AMvS5ovS1OsH8TQUpPum/KdF2SXaF8DWVmRRbtZpkj73mii7x6M2a
ayvRipIP6TMWS0qtVjDdSItpi5UD6PQtfvNSDkGKxIQ0md4piMdgmGqvZNnfC3as
6tNN1si3LIcPRYlhCR41kOuHWTgqzVfhKKCS7nbjYVKHJ1kpYWRM2mCT3Bv8gL2i
4Megq1ktePEYO5TqUdaJjKYWAP/IovPHpTZ4eCt9HpDhrt0LRkPIYnq7gt3EgiTt
FCi5Uuaal2YwXWLo/ADROKLyLRKamYPUjBxaGPa2CsyNYEQEqthTlpdr9LGjxBOb
gmLfQwp3MOsBOxP9FSPTwvekAPQEpE1l29eAmeLheTCVbWq0dxJuSp4ySmAfIg89
fUJBv9d4SZZnPb89h1ln9XoJWWzy3MgPXvEL9vkpjxrpfs3yrMrLPKYlIAWSAkAo
pTmrmyAkyqhpfVQO1rOiwnWd86ReUcMuTjUDATjYcC3kAp5E+zSyBkKw6ni3WOGz
6UCc/VnmONzIrBmCUwapMo5IjoqRIWrQNMSMeAv6Hf/MER5L6RgYuPmOQxIwxaYV
yu6d8jqy8BamXDoQdvhIFgCVbrkJjoFFNpPEKwUg1WON7rqAIlC8f2wICjR681xg
noIFSvYM3GzbBkc5poK/1Zb+C3COOXJkbDXH7woyzsPt/tiXIOA/IM8FgwoUGmWv
lY0AtAxJOwo4jgDTrwn1XM2g7oqvAmVU1UCLlyIBLm/wAQmW+hyPsXV0nf8rtMxh
UDRLuzlaO++3SfH7aD872jAfFZXgZ0ywsi5BZ5ARHrybF/TuSOWmVggFMBGYK63+
cXGgiqos5WvquUSEArrVdJeMkpRmQK3q6JPV0dG+pDT7dRNbH3N10URoDCXay/DV
egst48xqLbjQMGXmvcQPF/OdpiGHzRFCWZrsVuP/hYsb2nHYxM5AcnhIFXz4Jubt
3BUMH3sucQVMt9L9A4Jo/iWDLtqPAtcWAuS61Q6otmlz0S6OxFdIs5zh3PHKmpSO
fvmurC49/YSDOM9jZ4wAr+aqIyjTrWsakpE/8pG7N5EET3cQXYUlAHv4eqSZxNE8
tzPxBDeJW2jL76om976xwYj7WSTUMwhW9c7WuM/alSV1kd+dVVrqU4V520TQC3BF
IcBWhgkqDgeDM5jIqehSEfPGQbyvDbzfcmwgFeOHSVZrKwqWww3OIhkSk6DivM/o
uqbTXFhQA0ZFGjjPjhPq7t2IVBXm+qniW8Ejbtl4EZg0eujyCGhJxRym7RRxob1l
RVc+0A8d6ZHm0F1VYAcXfms1E6xcmm/dJZprWrc8vR5gFFe4QBZmezHCIhmaXnaD
L/yI+rjk8pC75cwMOA6os7heYPOIkwldxU1Lm/Ala8eYPNw9vqxCOZ3YmcIWVbow
olRjOvP1PmxNrYNyPRvd90ny6YmUoluo4x9O9wmcd+4msYK62Mmzk5DRLMsCd3tJ
XDq070lFst1BcJM+rMbRIIciuJ1pxzZ1eNNT2UEErsMKHI45Bo60ZmC7rSXRJSav
3Qqj0hb+kwynivaa2k+tbCwjwyPs/q7Zp7e1Ukrh8I06i/JkiN3rUkGRtQ2C8OAq
tzaLUx4vYdjA0EOzrARFRGyQOhfAcBrKWjGmbPw9IwkaoprjZsPvn/Uc/4strMrO
SQCwO0Y+PTkyBuyTHx72040/3L7UCi4JPfS3nxNbKQKGBXjOrjO1dbnJ+owNyn1l
dw1ixArLMOqPTq9a8L5gG8ffbyEgz53tLDCiyHunKRJ/jcMJ/d1voTuQKuO1k1GB
Qtu/ch9f1BLYmifSJxMmAX9fW/etc+8BaSpOnivvU4H7eAabCZOi7VJG2JEsT5pS
pTUUyMuG/raQM0d9xNCtMZghhzHUv4KYy/ZPMa1wemtT7IBLd86St1UnLd6Ty7Rb
to9QvD8IKh+73EOffwfUiBx5ZEP5CaLlEMPx18YCgbs9cA2q7sMe2GlJo+Xfa9Bg
wsHJhqhhCWQrG/sggtEEcEPz1u/mmDcoG06hG10PjD5bs2ZzsLOGyZW4oeMJNrsn
IFBkodDYPDtgLZfiFyRKl6i7SOaB9cVG5xr70SYXOjZTNNA4JapuTdCvA0kE92V7
P8ShROmLs3LsEuIdMyl4zp1X0jm8JTpWmwvSLMdVAZP+YEZPzNPS13OXmmi0XenY
KTCTvqlOlxi6mAs3vDJFbpApemaPpxJxk9tbK1oq0F8EGwjwyBpXGpLHjfTwTCfh
9e0avLhwG2F1A3GrIG0UaS3FQnxCuSB/vmyhpKg1xhtbTTgDv8V32XCrYCIpAAAp
BabG/mYChdPVpIS2W5P64mDOpSn6QJJZ7SoRZFiOW5D8G4CVq8qNTUfRKynwc5xR
MPvy3w6oiuMeURvemumhc86Ij+8WuQ7rbXThyxLCIiU3ffh3vFvcBhajMZnDBT0J
SF/PV8pKQnIO4zCVWMRSJPG94XcbVfYVLMIBtkbWkOtd03VS/qaqHMT6v2eckmrT
FBS+0ehvhKHDuWkU7p1uaeMf25b4hzKkFnecf7PJPWS09BJVB9KwgWyuYahqLZKk
QKo3A40yOFRjZmxl3fzuDPsdwDzb+V829eRQCT5DdSyENU27mlVGnjWJuqDx1z0N
Hu5a4JJcpBv7lUuHz4qic4IyaheFuYxFw8YN/McZ5LUxnCFROjY7eTbVTaXxt93x
MGi57yCWQScX8fNZdCNVMkFrLFY2UmsbHYY2t2nZhx9tsiPlskjPRTyD74XoB9Kf
MK24r0CxqvDZjXSt91/2IrjUN7LzDeqoKkZcP/1e2/in2d9t9VoxzXOq99FBbXAA
Sqv918sxHgs+ve6djduGXQ1L1S/1ksk6mGidD6NpF7BXkLFO65nFSlJqmzPpKT5p
O6bpncz0SPtBE1Fbf5loYJBvs/vrNQv1RTuub7zBG9CrzJZv8Ql5LM6yQRYTG2SU
wRafwIXlJBDG3IJuYUhwZEoTMA0EK67FulHZFyBBqmYc0GvQqEsW8hsQqLF9+KoD
rFo737EhsVConSQEqiATbr95Eu6648jbiBC6Bwj0nMim7Om7h5+IF/CHutJnonT2
ll2L5LSMdK3Y8owJOnLszoV/NvbsSv+XIlauog/E5qc5kMgdcEdAUrAdDYI8ChEP
NQaJpge8RD3rIwIBD4d6smASl7KuFVKktGJcMv+N4wRDQuXtEpcOXhUULF+mm3sj
iP129aMf3Yf+ePtRncc5MQ3MupCwZtbakaEcPIwvJnyShoxHj3Wnxc8w5viioOgQ
1ts9udxVwAla/+JmwZ1eM5Cu+FzM5XLMk+++bdj5LmuWzWK1xxMZeLsPAitAYEOm
SIChs8//pmIlTMqZ0ebJqxqdpbcMsx77Y/cY46+EIPtCewKFw9wmJJXj+Yqrpjeu
TncJrwZQidtgcy3scY5/8/bU86eZ9rpbt4KZPFg/2v6hAZxjHi+UwWrx593FRULy
WRJVVMAp4qfvmj81Hlc2oDGgSDhKaM7Vvr4LP7y6ZALMHmOdcWW/2blI5M5h03/S
skTJS7lvgc6RwxxZtzUWaJUfxiqA/hy0SrUf+oR6hORDSjdytUSRyMUg083tbQu9
gtgIKL/21RTKdu0d/gXhvJi6dwB/QtXt3Ca+0EhPOlBrbwnPuveugELISZ4ewEgo
Brsm2ORucnhWzJP+44Xzyn56vEgTqfQ2LHpy5k3CcSbYeZVPyqPUXOzEKI619Zqu
njA9X+i+/Cnqub+hufGb+b5s+hRFW2/MrnPc5RIPGcohcvHTaBsCyEjZqRBGflkS
WAlmcFS+6wDETHpUaZrmPANfoIVK0fVuKvF7EftjmLQw6kxialgNoF+Jj+uIg1yv
jdnVBrKsTV7GWPVofodBDTvzOnISxqxtr9xcXxaiVCjxo5FliCRUbaFlreOyxuFP
i80UVbuR9Gomo5dIEWqFmtGw8EuGd2Kh6o1EVILjbyrV9dol+E8dnNXm19EzSOIy
XQxn8mD/0wVwRuyUePo9bRzEeZrEjM8rrmVMOgdFcXYmR9h+hlwp4y4lXWQRH2LZ
9Ec9bDVFybInisHooT986kGa3CQiHDAD/QxsiDBzL7EA9/VoKdoZVzX9hKRaeygY
pNRMwfqNaGYwMxmY70xyl7rjaqrJVd0+ihkWmHZDsdVVETjxXD2TbwaoYgxnjHfI
GX2WcBT8CmVqMbl3zQNX8ObZ85T7a6DjB2FhMfQ3qpsDNtsrCZeDKkHRiGMiw443
PoyoIvbqti/TL1/ODJAc2QfmHWoNx3fwei69p6IrLTOx8RPWr27pXI9/TXHjs5nv
MS2ipJ1fqcC46v4J9IUUDR7WDxk+S31vAyRjnvXzSOAR1j/EXvkKeGHIYVsCZen7
CwpFgV6VgfTIIi5fFibI8E4+0yiAktGqQU0ig0oOBLszC76Q/d5I2RGEUIQ66t0X
/+xEOQmVvbj5OqTJ9eLGlIoF+RHvt8JyhmHlvpiPz/VTdryFJEVjhvQKq8w9s7/e
ttGUHcOzrgZ0KMG0b5ZuZFicnHNbNONlZHf4dyQ83dXFdhUrI9jXucs+Lt9Agxez
0WJcSHNCq30peldcj4FCl3zW6Gjbg0RkU29RWqRizMnld10b+U4LqXTmHQTpLDvU
z1li91k+ogy5AasyKUXZspe6qKPSBbdLBOVDdE4CetK+JV5hKJ8Stgduqd1GYfgm
F0W8nzAImukZjcYdj7h6hKgA6m45rtvucxWbnba3e9zcK5cznZ8fbfHBAsDWFxBP
WlY1euxdh5fYJoIOTCHOzWcrLi85q5JPXb9iMo/hXJWCGj8KZW07F2L6Ycgd9a1p
Y/L1o0fuSRhVUHIxvGOvAOpFCFrsE/ksVXTVsUMxPp5bK7IwJWrrZpAxV5qfC3BH
ZWH0PJZqAZxXZZWx6TvAJBdJ0HozsOc9OkAo9fSCvMvozfhaPreasDexuyh0pT4Y
BjW9KUcYSl1DQtMY0/CPBkaiI4HzdsOmegv0AzsqK4ts/Xg1WxVr14h5uLz2LdJa
GDrK+kBVkIE/rBNJnZ2b3VOEnECTwxafF9/e9jO4OFc83cvp5eGA7pzL/sTPp98m
cvdFGdrVEa/yBtKUb4OpxzV5s/S2S8e6ccNNOC49HUENHokQP8ot/fWwRfS8PdTV
4a5JluvtzsPpYo789z2OTFfRi3th8e+B5PRKMD1PslfAKmy2x1ziRKfOtymZ/BVw
YIcxK/fMPSaIQ+i+H5UtnQ3WxEM+ksk6LtsA6T6M0GY2qozInWCS+8gaLLfDaTFq
Cz2BGRj370uNg/UmycL/E7VvsfiGGrTvs9a+whoPY2iB9KCRqr9tAwdGY2O70gnV
ddQaqllfPnFiHYUhQAkRARVylHNWW+XPngcSgz3S5gdR7pqTudfyrgj/KMzmyn48
8CWFo8WBLsCLVWtF9+kZ1Fcz4O6oj5aCXyokge8YnefVu1SjUHzxJndwGEig92Sw
7+f4I7Cgq4xGpmv8fFvyjocNBr+upizfkte4pPYS5MxmOGxOrzO4NTgOfrx67kQu
G/ezBPSoDKUddomcIi1spY5e3drMRIyHXluSoJ7DxaHsWsnyneUVQE6cEH43G8U+
GfURhyk3cgcjxyGiaEc23eQvTpO0Yu69eJmy+EzAbJUMV4cV70t+M8oY2/87esE4
B2i9LSjjGd+LWpzzmz4lcrzyHM8VBMaewrE0xvLL/zq9itOvBiTU8SM9eltZSQKm
xWOu8xoiSdZeIlTW4H1+yyAvDDVeYECry0A2f0qOn/ELML61APubmji5jVIxm96L
wD5CBRuY4W2lsPoDYt1zOS8yBDwBZ7QV9WBFq6/SHRccu7Bnhviu3GKYGpiOKBQ/
YN4AO/BQgomHEBZXX5JJqYSsQXtvajb4M9WJu7z/du895f0rG0DrSo99P87oJA2O
ryA5nV/SegpLs7L8AbO8eO2qTEpJvrOG0PrduffKaYgpav5Z+xEG8mBdotC1cF9O
CrbRjzmCBXspcsLvLFIQ6qD9d71bA45HohiVfFNi09kdr7fmR45lexxteWdueHTH
EcgY41nvFTTcTmAHZv+/5YmrYXZTZ0l3jpot1EkjzQs+O34SEv3GE0CuK1XIHj4s
5GHfHaIjbT+QCK2Xmmc0yevp+cfcmMYBoSBVAUjVGO5qrteNb4MHPeQ8Ez3PlNDt
HQCFbPYT0vbvWm/fK4gtoT5RrzqVzL7GA6QEUYZnbbZ+PPoOZ7TgQ8x/qu9yJQHY
24u+sG+BZsZLVUakPyUw+fuLoa6nlG72eBsheprWfeEk7Act2UGx3csKTbB+sKjc
0u97uRu7PRhL2HqN2/Y28rX4jYz3k0KktmW/owg2s5pe55BiXd5MtndD6qkVCmOP
CRNA15qF82+UUS32NbntE8eqILMgPfldoDRvDyLhifzisN83uMCcxa57jy4Vdmpx
xZ3ZkhAPJA5AE2tvg1aQFuXlMpsOvtDXS6x34FMfkIkfJUNH5/2qPC2MH/AgMK3i
sK4/vWMReT68N1/Te6b1FJoD5YyxzkiWnH5OSKZvmmq5B/8rSkbEFGgq9VQm6vPX
txyH+I2vgYq+6RkM9fzMxQkONZZGDhpndh0SlD5IwJ+ma+PFoaRuKeiKQ0L5Cnas
8Z73wukYHA4I9V0dqx8a3UN+eSaxHtsXdL8c1iU4QjqZPNQFORRPBfZrE8FkIgKb
pKOina0jL8NlX9rfQZLWUhGqSZk3IygKL5Bo+Y/66uShrFiFl8I9uYuk6XjXBns7
1J8emoIrCJXhIm7HAPD34P6ZF9lMkATTRPp1ewx7sCrA0nw/6XaHLJtjq1SVsKyI
Xw0o0BPePDW05Si/v80AkwOfaYSZDvk2k5iW2aTmTtxi3QXwIGcxgq56XTbkx0BU
TjI5YxPdQzkUllbJkU0R1AZlnFaXhyMg2nxg1uzHKLDuOBAD/IptMBuyGJvmCkUK
Cw4BesavhfgiUVA4ceXePJK7h3GV5gGSgsszZ6ylu0aHp5EWtBa2lk0zQ2AauNws
w+FppAt4pDUwZ9YAAVPG/igcheVz6NjnN32Axi11v47zYVTL3QtGq8iYebgFxiTm
NiGY3W4V33V32orw+TkCAlNbg+34d6KPYGFaOm1a5G7RruhljRzu9zoT9sRLUVd9
AMsnvqE2oQccxGWmDytme+S35ZbQ8ato1ghY/dr+iH+0sV2VSXaE1xmqYMi6nCwz
QyZA9yxFmXMCZFHpLWdsteRnUcHafw4+FsrpbeSXcvDsMfRfqVFlNQ/6L7WU8JaN
CNDj2GPgBn8yQMw7j67aTKxLKZPBFs9h5uKkOEq0rHfGIlCWcFwKroauv89jL3Cw
SWNJUtU8WKVERdZkkscvYMpRlTfa2LdQ5zXco6RH/OQ13M3eZgkAF1ySjU9QXb1W
u4Si1FQOjdz63q8u0IsNbVUFgjsXJsE3+pPyYu0dju3nMtns2ChG/GVuMUsDZHo2
B1DvyQLStmkxmOvPqSLhF7IBV4xKadBj11Y9+ma8zrHG8GDeYB6d+VuifL1LObxv
cbDWWVDfPUa7/b3oYkexaXIRbAisjXjJpqZGk5J3lvAo99JwfiIaYASxrs/MoVJn
Or0ILrNk7aADJb59OlICJbFXxYXQEdM5zFqUANW2bGBkPRxIRqutZTYIqZKhR1K7
mnBfkI5ZVkLsmYw+7+H17R/BpX1LpGwUqND0JOF+hghFZ2wkRaZFfA9TBI7PiF/n
kFSb/CCfDqhSgrUxUs+T7xz/k1V0F9tSu9C0BxcHquubpmHLuGcQ+fRDlUzQyG1f
+Jicily2gLPSGebhGFtjxIUDHctvrix6z8jGiVa9dOOpmZIZTpS6JSxTmbgM6gQT
4ljBGk6Au8l04/r7NRtWzs8HsDDIyc23+PGR8/esidx/iwFwqESbbCBmL9xYQj1m
TEj+iuGWzbcbTyuLf1GdkFtwse6yoN3PJK+Tks9WNrI48OrljuVb2dcsJgLrD5Yt
Ax1Tvo8l8lo671xfNyNNTM2yRoUkv+gUt1AlZC9Z2uTdu1EfHC8QDy+tYN2F9boS
rPtq1HgJEpcrlGM6Iw5gKMvQVJZvQDVnhNeunZBWeoz/88U5cK8BE13uWVHy5xTz
JsMQxjaTla0iLtp5/GahmtZL9SkPm86d8eDddxcAlRO7O2IJlsAdm+pdIkJo7P8a
pJ1IA6dghJIDlQ2O76YOVrrqEsIEVXOe9foXNQaDaOPC+KhRV08+Ul5yd5pyeolt
ILtwdd6ecIXXkp9BNV9TZTBeSitqshuZ7AV6UCfLUHomZ6QHo/5YwmdYxmfAApO5
vME1blRmanKbsFd3ClTfPZzF4jNKgm0udR15hzARX+1bxZWjGsQxD9hJayHpnOHb
qSFsxKfDJqAdGWVRM4AhmVn8nhoH1BCHKWC7SRCtaKNjmYgLZXaIs+dSCtm4DwbM
/s9zRG0JcZZ8/tNHr4dn4fmTKQO83Rg7wDqRGkThfogZy2c8YXQ8fn7g7cKXTTYW
GBXzCoxC4KF2LjxEutLg/wWD7Ux3H4d1qGhUMi1pnZZVWmMBBaGMr5QQAwBHO4LO
2iAj4o6gtZmrGKbbhEZ55+LpDf5lifPcF9szJd3YWUGGyjmkeaovy5bhvm0ftFtb
x9YrQHiJz/7P2R8gdm4TXSM+5P0bChWCYXRm6ayZrcl1FInUYzuLPtYf9/xa1lun
2tfKQ/n/NASziaKytzkUpziT1SwrVX5DeWW3pCKRlB098vMeP3DD+ZpyTkl1V6/z
6QGPPbJ6N8TU3QHhJ8eW0re6JgkV3gluvy9AOCcPOT4mmJeA7jfCbtDpU5geUHTb
48GJ8AB4FuHSRZI0zP4/qvbuliU56H+Bsx310RAj5XEuRkAMeZsEKJzc/9kTAibc
EhD0pkHNbqP2RioUqDOE+/i/HLgO9fObWSNwNdilWt5iV+rkMAuj2gt5V0BaulWb
SA16nQ3WJS8gV9V/czdHrgedoCizEFBv+fbA+3moQcYDknX4NvAZ4ljO7zc9xW8m
wZ4tXeD8py9eDcDjXVVqh7mQ0bQy3aco3wcy8J2kZdLzO8rB8KLI+8aYjM3kBysT
kpOZz5j8e0CAK03FDlwsBBxm9s711sHrLgkdJTHB5TO/jEZPkbjpiNwFd3Dwx0sS
gQwtbfcrbjj4HN8sjidW3sLv7mgqgtA9ZR5D+Nf7oUcpgpo9uVyipFOQIJyUsgnj
EZLHA4v0avBFfazKDN3KqcaX58IzhkuvsQt2GiCXNW3p4GZRYWZses1FyuXsQRWO
qwSFiMUl9Ps6rVgO2rycngCvUBZC9WbI+hEXylXOr47DTlFuCNSN5a96AKLpKiFz
vvo2+k0YDBQMRHjdyEEeRhy4wb3rKELmttW3ppdXCa5N3bdhXpQZy5Xha0cSm52o
MA1pm43z/LjwjzznOrGjxmmUW+LpoTiEzZxcyx9v9Yb+HqzOh9cpRXwMvU3Y1Bge
A6dWwiUPE3eLLdR0DrU70soeXsyLGDedAuBtOlDXbRizN7U0zjYAKDgsOsYwNt31
7cgN3JCDyN6HMzQmR9QVmsjwyfpflgXVnmLbnv2xUAfsrq0SXXT7Npeq2n3qafMk
E04IpmHxQ43mbKe6uWP/q7hLNCbO5oMPtHRlec5lPuryi1Z08tLxLcqaxjNUY/jR
2iUsNI0SuG0yVCRYnrl5+DTB3WnVlhncm4gawd26mLqiTRTiZ9LlNKx52nIGO2aU
UFL06NZEw0OP38tX/8CqAFEby78CQ0GcRRtnq8Wxo5sc9eTa0iv/NXou4EmNZ4QX
GSS6EK6WFhTzG3YePLD0KY/drvJHZp27KmDUowYCPRjqv5H0PvDBMI3t4rZVVYFT
nZdAc6u3y4IE1y3RvnK7MXaXYwWwM1PwhhBmKPwnb46B9AWuHhx9BpiecMLZpl2m
oeg1LUip7wBp4bqr8VH9dBo/9hDZxaVlg5Jgssk4Zg8PvjfV4H16KdXzjKFpxq3u
tduIl9/rEfs1yiPR1am66TuQbKVa7BlWeeOcweNY/1LDttWUTD8u5u9vzle9PBZb
0FyrraUCKTRztH4l0wEHb4mkDfQ/E7kPRQwtvaxuUuCCbuM65GAURItAaTkDTe4M
+ezvY0M/ykY9RMxG0rOI4KaSxeLyr0wkprax8WVtp0ML/dWXrbZ6LMiQqw5sCFQu
BrgaIIRBEzKXuumA2ep2EbqyMjuXowMLW16ztN8y20Z/snhKnDbR5y6qQsgog4D9
wbM98ZJX1/RP/oSvNu+X0c2crBU9Ik8j8gsbRCiEfClGvuMM4LmiaGgXcni7kcsn
JPA5ni+AhEfHlSSGw2EcjdlxUYtrS5MBFTqLvZ5KyDs8kqrS4OL761lKIQ5KlBWD
zQp42Eo1tn59LMTa70QpWte6I6UfKhHUlV6kXnPHo6akNLuyvwcNQ1GnLF6+3otH
pgr0M6PZoBNMfA8WmHACCsUs5FBtBxdp7nK8aGHfoXM1yb8oNQPlpceXHa+xIa7d
kAAphTeGOIW90Kup8Yx1Gkj7V3xCrf5ejnaXYuL2wtj3MGMmPKvvqNLbrhG0TV7u
XeVVOOfJtTouMhOSbaq3bdFM/5oOcEBLSF7YjZqgedW/WjyJhdYwKCVjN7Zl5Rc4
WC4VbbDzvm6gboPkKQ2G+XM92FpgSXgHWHKr5luy4sSV+3JHTmzD5PJ2afmRaIrA
15XBFqZs73lIKJDBneOkTHp8BjAe3xQuxrFR3/Ne1r6Eh/vNAN4wOSszd5ceCK+N
JdDfIaiRGTiFHKaKOVpcJmxVebzfhypDWStKrptlYM3HA83Qn88IqypvvhAFt987
vheDHiTviBjlcQ8BJypIq2AU65ctw40EVyY6KY7gnUyOJLhiXYCYGJy2izEopWZQ
6xMoMBmJ3pqMrUlaj6gsc9LFLnslhnW+1P+Hmq46Wo+PwX1SHUOS+o6R5or2P3pO
ziXqwOEvnYiIYPoKBQdLDyYl8I303phM6ZPpkeKw5KlQCpr3QFtp+XoCrw34GuT2
Bq3oGROIIeH+osudQ4DsQRG+cj8UOD8g6ZWLfNfuFCIfyp5VilLhcJ8L7qprMO9h
g3HzkwTw+XfZEmSE4M+SY7quaS5UYkawSxTkefiiGZ+pibOHrPBe1hB4HcGjQ24q
IFp1ZE8nvZdGnmco+UvqaZOYZi7sAfsTfLM0KMMHBW2WJt9SRAd9gL7oanemPbGO
tQgopSjAfAIUuMVmcrVJRxe7w+6DbQ5hcidkclYIcsOaESp+iUDhFAn2dTZBsZjP
/Ed/kbFitwlyYU+/isy1f3rBsGc0qYoZq5i0t1JKmZ9/U7lCM44qiD2+PxveA17l
1z6qmy9rFEVxqcL5lIyzFkpQ4R7DeVxFbAJ8zG2mlQZWHTQ3VV9JbE8S8e/TLuR5
52+cKAEaHOqzXvoklf7Np/UZUVmNPbYHTg59QCtSgM1sJFnKAppvZJi5nmrwTlJn
DZ3nyHoZkULozb0CIUZJ/+xub7eumvkwt/KldiZP64Yk5EUJTwjLIVLSzBWRSWEv
Kvvc/kpyO4eEMRdWwdYRPXIFIri5/WasC32+pvXACuv/q4c16+Ma8NjTw9Lyj9Gd
F0UUjWuJsL/cKF19DAqjg0IoMbzvfqriQrQbVXwqRPmzZMhPCEMTiaYENDQvxUO3
ZbDHMp3DaXC0tE5qUkDebA37A0adoMOWR7FOp1/S/c6Amzbs/NkFKxMdct7emjx0
BpHH0ERYA4u0TSpJ1ckHwJsmCCnaVNZ8NLusSHwsBHV+VMAkSGLNn3i1IIU19qps
Pm3cxaB9ok4oDzE7znSKYqi5Q3QqWHCHg2NzpuMnLO35E6Ud8CbDV6tLRJvfF61v
cpkMSGFvqlTRThqdK77ofenaco9WWFEMOeIcwwjE9H2gJlvmk2ZaUoNSUQNJTz86
N7uqoiomQiPEXHqJ99uUGvCrFz3RCDE8d5GSgMABt5/7nLiYf8c0tp8vSQSavGvV
hnFwFhWZHTFpV85GMMiJ7KxHlwrWG7UniL01nnB6FKg//Gf8K0vJpPNtGwc5cSgB
ZLoWgDovzK5rzYyqNtEgNyzToRds4ouz4r91pQU9Ln6egclnj+fLy2Imv41qPivM
Zklb6EUfiYqcA68KBKFU+Ee01DqGVKToxrDUHxyAVbLmz9Q69MJ/3APENeM3PUhW
dERJinLMuNuMOTAA8TCMSjZzl3HNTCYdJF0U0IwIxIFWWcavPeXRRId8BuUbzfM2
/auYjg0fZg7wrnXlF2V6Wql6UPNSbSri/zjAsoERXgX0fzYTmzPUuxeWYZ7MncRn
D6IK9R2KN7ic5RyEW2DdVDX9ZXtfOm0kFdDd070GyyZ8DpOL6chljeT5uaToIKk4
j6dXHW91ZH2Ht5k5zXtNiKd8v79lIIBFtkcwgMTdgkYEtqW9XS1E/V6VDd9q3FmM
MF3to0hWVK2MFpzeDwYEpAdnx3V/6hFz4IdYGDURkFgFA29C2MYs3n+JpjG0CUva
Sk0u8nJ3VHTTq2KI9VS6jSCM3bWgB6Q86Ui941JqIKkKGlTZAIJIjrAnmDTqQJ5h
CQxobiF3KLJbW+fVoAPMhA9R9MuuQattJqifdw3s8LXdBLCs16AEsfOpNdVVRxRd
OYNPHP+xWA7FE4H9zdatHcLyYtTJB4SYbRYF30knu2LKetbuQZgdE32laaBE8r0Z
Ogr3zIRunigMdssuHLXvWLJAhQKDHze/HvSJY4tf1gg7P6tQvl3QqFL2ta0XQ5NZ
kiFdhsDsuy6b9ePUno4eLcEB/cYVmURZuFe4eEsMuzqFY2m5m8XXcvPNNUeRh7es
mHSuOu9pz9Z3OwpUkMQXjgsLc6OA2hu3gkjENTrL/1TpEhik07X1BBvvwbxCeYgP
RCnQBdeMXZ2UlKkicNN2VvhckcsqMT/RmP1nsWLNo/gV+niMgsURZKXQtAL4e9wc
oTWoJ2+i8Qi+A/RSuk+YCb/7kKGZno+PZOz/6sgl/eg3sJChlmctsDdotaO14HEu
qp7vvgH558WUIK58qxYAECCrXRs6hTD0x2wFXslrxX0Ca/q4wvA571keYrTdI3NE
MrkuQ9W7PISOecGbO2zH9CfUj9su71iXtoB/4dUbIU14l4trKXL4UfAL/18p3Q2B
xRa5mgn67Z+US5hAh1aHL0aJm0ImpRnXop6tJGKp+ci8BvHg4U2q/pgYEfGiaezQ
DpEaZdazy04oK6AO9R2QupL4Y9R0NwztWQd9QzMErLT9+Tkdb4Tgd3WsQXjeB2J4
wd1nbAdsfy5NSWIHdVLb3ARQGHm17OVpLa0C585XJ2/yXwHwnueA9V0f1Oa2ie7X
IIu+XRLjFoZioojhzqptGo4wweyvKSZP8k3kjqygqIccqMrs5rgFlLDOQJasVowE
nPXz/Ai+n4alol+TOMmN/A5W8EFwsDQAyPXxwBAq7wepZvpxtj8F7sNFp1UsuJCA
DIFYiF0nFOa3WiQBvNCSoIiFndtFm3SaDzLfC064f5gXQGGuJNrInafjn+fLT5MH
s6HKXEvarBzEuvQMZIgUBq+iDJKikTVCit4DvYjGy1QoT0EcEQ98WwnvEKcvpzOW
xWeQau/i+q6mYUU9dZX2lk9efhHz7UoDK5nXWeyLn2JofgtZMT+ktvL1AZjbPq/4
FMBqtihvAJ9HUL6g4s2O4PqE2Fm8elg272WGJHM91dV0AyDx4S9nb1rOEiPHsWUX
rd71deJ7q/tYY72mLGl+fQqt9GpTEiDPiL38oFiTMxyAQaa6z2CHXxtq3NkLXrnK
6ROJWPQe+Pg8MnNA5AzRA1r9VWmKkMN1eY0AKwqV1bN4ShehWGP3YCvLKt7dvvq9
ortxrRsJJfEg03oQWtcCwwiaD+4tL7RmQ/4fk2DDeSmAwvlXj11iSr7lq/oFMmp1
KvOVaFTpxFmVsJxWTxBjiPdtJcjFTHKkUe2u0JH9a0NaCYUwIbXmC2EnRUOQib+d
9fsUC0En50EjS2SQLTo6EjQLt/8j+BMM+PJ+s42+aUDhu8wcwPIO8itAwcmaoU50
b8Yh2janTgZrQ+n7ZNJKHB4TaypZCoLNRK6YKmpdNgBqdyvbaUMDPfXXfi0Iia58
M2LEJyLQ5fAo/83hdviD6Wc1gkrvPsKi1PX0d60zFwgRDbG7P2KV0XeLvCeADxBU
KFPVzbw0mxA34tA3IsLUU1bgcR8FmENFSeBF4dUjaHu4Y4c0qjHbl7zqudAY4YyZ
c6MPLXreZRvzAfXCa+2V1syBJHY/sQLxy57QArLdUl5dznzBkHchXUGUnr22o+Qn
uczseNp31OCk06pM1OyzZnJGIJzReyFME+BQyasSOT+aEstyKPcPFuDKHOUNAq/a
9SFOpIsmCY0B+J5ElP9wVmzN3fzKMLUmh3aNMT4DhMARH9u2+COFjtx+SkuAF2zb
wEL46d/9YJijqpnqT6UqwTVqrmsuFR8apmGTZqFxMJPWK+Et0i2KmdnT9fk2iJ3r
8MGt1lb//FdXIuWcbtaWzicIea4kv5gcthkZXKCIzw3UiXq3U8tPa8VZ2HT4E7oU
ulKDlZe8BbG1td1T6ebzvQbycHeCof6A8tKGTZvCZ2fgX95ecLMQMDQRslJxDkWI
m0MaNbgYno0T3X+ppOTzpJ/oCASFjZlGKfGDtZtXZzQjnOc/XVjJv8VSTMAKWYAt
0IjXJFho/x/wN/lyVy5kfha69mlTGt6eNQfxlKBA/fkkEhqtRlylMVeNb7wm70DJ
wZPF9C8zwdW5C1l4DbqW9SbW59dYpSWsi1FjC+DGWJk1SD9msfIimJSZ2haYFnU+
PHcLa+rmyB7kUfI+3H4REnK9iGGwLHzrcCgt+WTPKF8pvTsgpD9cV8kfuFtq76Hc
L2cnFJ+RotNXxaX38/G/VOP9DKeo6uoFULVLI8l1cuXR6n6jiHXNSRBr1SfmhDl9
RueQeB3J12m4l/h6hTWXBn5Vezw62hDpuiUHMppIWShaQX1oGx/kEDUn15Y025Ea
I33gqghSNrdE+IKBguCBvWlXvftxefCHQ5i1PCSGKyPDUhB0oREpXq0mt9zAucCh
71JRmOJRy6UaCtPFIJkRa4pUqjH2/x6vVhhrT8z03/Uco/Pxm65NdcNR1kug4Ff3
ZZuai0DHWsmYe/ha4nYHv4qbVOwwujTrX0osBeNPjyq3AyPnnQSqjsh9D9i9WJ4n
aLrs55+lIo7g97kvs5CTpTel9F231/+dhLnRmaNjbG4SdhaJGmaJZdW2/mBn4FyE
N0jK/6oaY52P/A+RuFqbTk9Q/+FHIFPrBRzZeUvhRWbVlfFSROd4kPaC6Xdzq99A
EILTq0AO/7N+0tlefjoUlXJRwycr9kstXKHdk7bLlbj+bIrhTiI1NVgMTTqivfrd
Sh9bSzd3JmgpDWBvDDXyCbsr6+ZwIX647MHAgo10XTyWLcaLQyt24/r038Eualbv
on/HSxCRX6uborFv1tI4Xs20EpOiUt8PimeafOBHz+X6wD8q/KO2VN//53fXg/UF
p/xIOfklCYEWLRVPf8L7XkqnllDK8XBaGFM7yOQ4tBjtbZ3VVVQujIwEATp4xfZe
tqpCshYYTnOXa5P7qyRhQ90iAco5525GzVoN1HWsuvIra97HoEUwp5Uohqxqh/l/
CeD4fjk2UqG5lp93gf427YQHGxMISyMX2RvWl4mi1H9hOb2dYeW2d1v36wRTJwZF
7eNYf7fjfGxBmYejPvLGIdlYfnDma49VCcuqI3zf6rOxyfbNAXanCE7WNCEJHMHC
pa4S0AYXlLsWvxpGw9cIKIKfHHyoG/P8N0HAHMHfgEnizdMOJh7RUa69jCQHxIT9
ntLR4vC4Z/U/RMQ2GNqo1tgHCTa43Osvvpcon0BdGpnPEkwGxJe8bi3tfC2b+2+9
YyieoIZA2QELjpdlBB3/vVM9WOT48xZjRDoChRgNFBPdAymzlx65lCn3M8BegkGD
DLkU8udFBB7esyn5nHTaMznZslodhXhUTF1eXIgo48T3SCamNCnTNpww8q0Neutl
p1Dc3MgXCr6F1gpgfaqYBHg6MRtIly0b7orkaNv1AzwKFiBBEgR+/Z6t8UHBq9ec
oMuiqgtAS/x9ZWqZm2t/iZHN1hNGt9j0p3J3zSAsX2oqA8lGnr+R5lN4VjXeYIJp
gQcJLlS6INtavSwLh4B31T7xpS106w3frV83kCdaaN2sCH79Fc8J1meQOdWgmDNE
RDPlci7FP9yjX6izmVldkQ7pVDQ6Gbl2RYQasFThaNetsf3F+9MP9da81tcCoeiK
e5xw3jDtQrPEMfeZvATKfj6DAPLFFZReVcy1/bC//pEJbJlvBo2Qo+xz1tOjiLdy
fBSeuRrFT+lvFFVBj+QwGvQmmM0yQWGnQT5BsoO2gB0pN+kgz3jrYtC0ThvMUFx/
eAkJXmBNVCShoDwxXvAlgyXlVGOCP/Guw3nhxzu+N9vI7zW94ydOicIOunTXCeX/
4GBIxwD5oi0ZliR6Ciz0rXy/M6u2zDCElsVN4kJ2XyJB+W50GxU1DzZvL7lAx90j
J2K1JSbcSQtUBHHVdsAtajAsV1LAEBBiTlwgVtv9pZyvDC4xVF6D74iPC2NFqS8J
rYrbL3Fn1wwtlOxg5qs3enfed8G6C8SZtP2g7KOwV2NVJncOEO+sC34Jg3JqJS6n
Y9+s+eol4G9vODzQmpd88H7fLgIIUXzDO1ddCd/yX0oFaGKQc/h6RlbGiMuNe68L
fWjzFZst9LGaEb7Zstzeh0qCFtgtoKR1KI5jPpWoLuk5CFE33FonvwSYtEBUGgKl
nUANnfgjXmmbFivAFzfeyIk2PNNDrYRqBObAE3KBpx8akD6k7kKBNNlJYBwUTLzs
j1ip5ncdcZhk6XN3hRwITkupm4jWl2bo5+zDE7ZydDRwf4JdTNaig/29cJNEBBGA
d/m/XNwrgrzUhOYC7kvPiRmI2Rb5z1ipv9Z13jYQTC1297EN3di6t5B/k180hdwP
vKO+bKpHS6Rcg5F1KBrmE2hiRrpBIKqzj7Ja9v+mxWOl1ckGY/+YMfpT9pCFxv2X
N5FPufqw3orh2RDY1U/kIzZ7DGodJ7p7K+aUL/5JH8H+ZFvbxr6PwzSlWJaNYEHS
YUvWqviOd07XoVKnZ3nZ07Qgo8JTtG6WoLhGJBiLybjyib39HhX6xgfuwBBRuMSZ
+k8BEhzDf0uoYNCIMF8QrdVLrR8daoe46DpNzKHMWsr0sDtzvl/tNgcecDXdKGTd
h90tpulM2M9X/gJgwf+2zOTE6F87w41xoGsC5MdBpdi7uIq+EuQAxcBjceGwHvXW
mIsI3JFXABfr971yHOg8infB8IQ31EglQpZYjmyOfYJkzZcWEpb7wrimMFPTDk1Y
DyhOnqOrqVG95b4JHoIAZXY8z0J1+h+gZj9siaqKVXGQnZ8rKBAfALRLa6CaLzpQ
BQ/nWjfKvqma3eAGteFLg3qmM+Tc2sy7aoI0Rtmz/Wd6UDYBAp+5YWIc2meRIIiG
oiKp8L/6KjI7i2aI2UgsTaq69fpOGLpaU088XVB2C16qNoeyGkxsWKU9E2EzAYLp
2+iKJBnFhQtiEJMizM1FORsQItASNKEumiMBPVmZIpm7tGI8IC8CIjvSwOk/bWrK
x/xDoX9ej0T45GrOIUExgsgos+esiVANaLTzPgdgpxTRQ4U8SsjESShL8KE4XdbL
OkpRmJeUR/nhFew1nmVJ9X+llvG9JvaILSEP8OlMyIYxymRKPwmmvqA86Wfm8GRc
sToJIc4aJpOwnCNrFklCHeOqztkKzIO6mTujJ2bJtqKNeNw7mlcftDNuMI0HUsoT
DQJvzfpr2b1u72f9VnPOWWzNpor+UM1Z24kubsFoMWtmlUnjA5JnDM3ky8DbT/Dq
oo60/Cj3FJaE0uTBODOAGfDTyi2wo7A7ujRi1/Cz3w6+ypBBH/0lapxzNSsf7CJf
tvC7mn8rnmF3G3S+xfQ+L9el44fCcBAHD3OXMojLsXQWOhrign9curuA2Hh1VPPW
fVdmXm4aETDkLirq6lCZe/e/aGpS0wk78ndopedXOw9WBnavOw9XJtSW+mfQidd+
5CpYKpR32SINMGCCpGn916VkSytg7Nlmd9BXCfuEC1bB9GK7UM0yTGTS/pgutEt9
YxLTTgbn4QP7g8/v+p8GQ2aB1okZ7VsaVrXJMWGOocjlZNLt9VSyzUIZ9suPayhF
7xgQ0p+LFn2cONIHf6MUrRrK5cq/YBEexe1xIfAn39PhyS2f6qMiI+z626X+2nLF
rfjLFztRFnu1Cstr2KM9HqDEKGJMlbPtQ5jRlvCQUdSFZv+G32gVgBKsVRfaAzrz
/dRc/0OQWONLo7E21Oc6GHZhZOjxxPB4CZ5tgSHdmCYajD9yHExoRJylIAqi90fN
YVoLbOIoyvW0j5vGnVBGP4GV7iza/OkuHHQkbSfeFDs9sTaUR2bw4NjZFC38+3gT
5xKk+IpmrGPDiJ1N5IPz3RJ3kghiZ+AALMh/LlynxbdjoeuakrSdDfK4KRX6pm7e
Rbj77gUb/W2cv1RzyDgFA2EfEuC5XnCjPy57UJ2RXNAn9DxVGURpJD2idTqny8AJ
DciYfSIogdVrIyFtXzYJr2inffh3TrhE3mvKv3oMvPC71TbiFoaGxZwQlP495m3Y
ok5b/1kiGzQhpN+uSsYx28A+BVVR4uU6IbHacdxnrX9ADOp32SEKzVX7OfdinNLc
LCHmQKrleNcCXvKsQovqjl2bUV9J2kuJn8T4Ek6I4y4o20KrrGMrruPZnvgdSsL2
Qvv35j4AEQuFefnL2kw+Fhy+2QxbhHOl/+dhVq9yfzdhrYxXFmiDbHOX5lobI2YE
Z4A97VkhoRAsn20ElgcD4Zfuc+Tp+HvbGiDirMwfuhExo7RZod/M7ng2lPHDE6qS
AUr/535u2JkH/imqPQ+R4wcqUoaP6eTxOfxiWPs8fBaF8F6dXJbA4oacBgFkom/o
TjM6pXR32LvXIV8J6xJ2IUSyt3xoklm26QP0IOrMI4aHT63C77BrRQSR9kTnFJLs
ZbYjY2IHBv4hLMmAwwxKNp1t0BLy+qoT7j6vfSM6Cm55WZGd9q7MM4dorOtsnYzn
xlC30VJ6Cm08kAFDufZpNb/EPMFLyADeRf6kl+zCD5wfGoIFDM0xCNLNws8p0RZ4
BSfZxti3icbQv4j5k/1fRqjigCWGY1Q8lUuEJB/K1dw26TqdAyNajboHnY4mPnIz
W6589CXJLI1Ji8xXQPdA3U5UMHE0d/BmjHux4o/2R0KsyOlHIVtmzaCkMOrLNf+8
dc52Pj76lruNNxN1S0ymxVGQy72Em8V0lpIjp6Kte0R510v/5l+GPHzrE6NfmA8K
QO+SbBYC9vN9LkdbNf4MHMYo6C/3MIfB3nEno8uI//dUVean9IINgt8YGGJUaKpE
E05oOTWg+w56XXa2cUL0qzXToXzF0qb/Y9WxZ8IdeyvRv/uwSZPLlfj38riWW0Dj
qkiBbK3bNmz7on2n2m+/SU+MXwcpr/n8ITqGAqN8lGP/CiA1njUNjtSwxF0fL7uy
t+ISxCkKKlaO0gHJ6xbVTXxQaFx17Dr3F9tTeP1oUvg9lXYe8CWi9QK1KVRa/KaL
wwzseJTuilI5x2EOAkyoZ4cVTbFy0g4niaTJ7R70+hgjYjqNXLeBe4R7shcNABq6
yf51vGTrG1n04WNTro63wmfySfPNs2t3RqeMUj9rLuqYLv8hLN3Lq4qTrJf6T+ct
Hoiesz1QlyHIUrbLfYwbPINZmqr+/shuPh2nGL2NgCrt6kH9ImCWOT0fZMO/dqTk
gpNk6k/3qi/nNIf3SsF1kErE6PvzDJVIR+jns/FUX9ZdNk9Ks8VVgffe6H/enZyt
NAESjC4bbrAL4YDN1iR6nhDnwLjLV8GnofdHTPihKxvxiB0LxvNHbkYitRM18wty
+xOsaEe469ewEQctyzdVatr7DLq0iu/wJxBpa5qQcyfoW1MOytmyIr7ryxyiLc0R
xaylhZD7ryFfloiYksoNDLlZZLzRlguyF+7SniI0+Ql52sIao3Fwpz60HG7Q//yW
sHpSQ59ihvRbQTjf1ICudba6dZDFdGY+dxaFZ8muWjl/y8cXnx+WvZ4z9285Q/SK
wjVEEG9LSRTIKjsObSJgRpJN5T17NK5Mr+s683UNA7i3ZAimZOT3+8gMHFX1WDGm
bOdr+t36807oGGwehQ2S6XUAPd2J7WJ3W6LzjWaUA/pB1+h4Wsg4AeVfbwtC5sAk
DGucXf+mP6nZLEwov6g6W6wz+y6wbGMeC4WOwtO8cZR2NfI4X9lv8z/CkRdgVkji
NcBKgY3sUAdhp9/nQyb8MzntX9OLQOIwiZTcn/MUlt19V28vB8XxYo1zC+bWS7iv
i10u0Kwg4iuBCxISCBNu+EGFw36n/Spa7wpAf/riEFxmwSLXrBKu/8yCRhTc7DKf
CqwYtdQTg1A1k/ChDTH+/dqjZHHbJEUiuvzacAzRsncpsH3n3Xbne+Lo6WVlpc5C
yKzeHQjQvfJrGfLfXojfpxoZnyNlDqFrRkF5oWN7EtHcD9DrZOGFlExGc+DEIZCm
C8ZkDfZ+vmLmoUhT20vLPD3MOLhVot7xZFuIbExUwMM8T5ytdFNONB6MbFcJnM/N
2omnC+pH32nNW63xr9xrn1FCsM3MIqf8hh8OMsI5br4KU/q6bIOBnC9Uy06JI+XR
QGirNz295DJ3BA2mD4b+NB8P6jcU7DDPQiXPd6LJyaT4KNWmNFRV6vzScIuw8hE/
8yXnsATxnbdvUtb9CAo1S8o0771ADlKCi/IChZQkbLI+FLTQAmIelk4OJBKvjWK9
6rwKAmIKq4wnzdQ8DmCMn+/Lm5DBAr99S7Ij3eX2PMhknKzeT2r7YNRGVSeimYkI
dANWvgjourUXAVdzX6AaZHjTzt5A0PWVzZVkwtTTcHKRMLdT5jB0e+8pYhWbtxKK
vvH/OxdfsvGVHJPMwSWm1xVC6awJo0DLbVHbUSukigFEk6DLBTer5zRNjUJ5GUAk
WX/fXmgC8/EoNOnCDfNGd0A0lgjoFbcb04NyWrCQaLykJ/hbdFyGwOUqjhqB6En1
bZgsM9x7gTiTL8QZFrbOsK0vrIVXmq3uN6kAYI4Ze4zNDZeEvA2BKxEN6BbxJfwJ
KiZ+LEKehDP7WPqQXw+MGzKGCytIy6ZPdskLgf1N5v9IzOIwzHsLYuaeWxMPLxbF
EwNGhHRq63Oy6sUtNleDyfkSO0k/kqfLYMlJ/+jOWczn6jVorR8M9XnHShi4XYuw
WEMJrNA6636wDfpMxAGELu+nTw9z2Bo/OeBpEoqUBkjLOEjmZQqilH3HbwNM5EHR
eb2zspVYyUYJ6Kew6c5TVhd8thOwG7UCeasBokVDkEvYRq6RYRIciaTzRy73M7a/
voiWHfpn4ff1cEjGIC7dWKWHcaF0mufR53kEcFixVxJog1md0RWfQVAKe+W/oOO6
ueRqoqMae55WMO9neMuqGFLeR8BV7trA4acNADCOmsQjlwapmXl3Qu2w7IhKW4E5
QZGwWAzepO5A6XG/+TH1/y17VPEiNC1xh3IWO12+hJwd5t53dd9o92Wp8DIyyHy3
/DHg+y2BS+K9oE4UyttOTV2lalKb8yVwNNPvk6m2azPvbME3Awt5XTyIwMef03Zg
1iDosscvnqmKV8qp7AXob+fWNq8zM2f411RWctTGmhRn0qoqtUoV32y2Iy4L8HoR
xul2JcGr+RpQbfluyyWyYVrRvQoLDEeLLrcSGG6RAEOmQ4g2IQ6pn+zrLfZv48s4
O209eHcCChvDuoulwIIgi1JZ5TQv68P2QJh18opGZu5+ls65p6Bog6S7xRIKnvCm
UYngDCTElF0cU/ZbNqko8+cmabTqZqCgQmQgi5RWIGVT17hsxd9iUlj1u+tfqrS9
WCniqseucz+3CpXjc2XWTB3aBTN4KsqWFECvFjoSETX5owtHRV5QR7v8pFOTNgBb
SnpqRPT2QByxO1P0O92xhrKRz9bl2w3hzZWr1mUlYjidpzwLWdUFj6py4BkOUeoW
h5sXZ73QteHxHDcFfyPTbBWtUn6johrX4b3LQLe9zClLO5mWTkxX0UqB2hfIfQpR
P8dRwNemT8zKLwmt5h0jdMHauCpUg/LMQ6pP1L7HXIHqxOx3TLKpDL4EcEGtFBix
zJJB9bAHXohhCZlU6s81SRnU4tBLbYjFRd7yIwHjY/JIaMKVEP7NUpeoVXuRn+iJ
FsgbBPTRyEpIJa+59eaKZxcyZX8Qz/JEc7UZvNpIrdgonT5IpGvQVbyFY/m8xgY4
5ioGHrOp1DOJuPCUGM0eAYJ6eCcMYke2EjWjSudKh5Xo/2SXF/xw8vFvs9XASoU6
X7FVcMOjUJTD3FQSyXrsoC0mbXPOh1hcq2VX3sy42d2xMXgkEJGeDwKOcY23agoF
62nISIsvi4z5aG7h+ngKgymHzIxpjShqCrQth/qECAGpUOaYVsamKYMj7GOIrMem
8dcW4J73U61X6P9+MOeO79thrDu8En9JLwkfyHpWqPH8sPRJe0gIcrnph+WBvLtl
j/eGexJVzzDaynCZcR48hL1RNzj6n+CaFnUCHc9pd/VcBQjU8fYAHVmLH+6n+Rg3
9QBFOSuoRyADKgEBnGV7kU8qj4HbO7tn5dwoFSl9vW2xeiBOjX/MgKnM0QXjkdU4
ZsmpSCCMasQNY2MY9dcuWIfyeKqhB+xRk82bxUenx5Xkhae1W7KY8sUFmEb0qayc
B6MkcylU1jjMa+7klK5O26tRskEJtoeApVhRskHv+YmQezVN46X9XsK5tuthhG6z
t9lYuxucI+hdtSUkG17+GDm1QZKiWnura/NYR2McegHDxllkerwHfN32rpU/cNVS
7e43yNy7PPBPpnoS/95yRjgWvud/cSvj/dbpbsX/P4nvMY+sPewL28MKuhYSYWYw
pxSQVjZAZcj0LQCbaVugyqPtScGPkjBwhf+0XwrIM1pMSmCQ+P6ZxxI7We8WSsmh
EkZ0s0Z1XMZzzWBY0B3ox9PwbO3oDybDm2rWUhQ7SDHoTCvce/Zmsm6Y4xrtVCj5
YAEzng7An+X5s0dfmAqaNHV08LwoyGnEEBZhvh00+PpchDaZPSZwL00RK6WHJKVq
GU9BnfpH6B9Dj3kXOcgOW3Q6JCFfayt5iyb2vvqUIAv8ox+aOLeogAirkl8RGd9H
lIj35Hwhl7tPfQhecKGLmKvafcNBqIcAgfATppLAsJtDjyg/G2zECWuSr8IZtyvT
DGMlJU3+GFR+khmYLlGyrxfW1hyuH+enuTCKmzwWgJgkhhP97GZ+068WEDsVY9A+
yp+rUHsC4Oqc1JsQeRbq075PCGMOUTl7rHmkIAUuh0XUioj8ht4ivL3yZe+QlChe
NXB/7uyhCaAnCriEalLLTsC8JIUyMIyaumeP5HagEreCYcJoMJklQN8tWYPKJ201
MoYLZrENeQ2EMmbjYwOOT8VJF4ixmUKVM954a1WOXiHM/v8HaFT4w5VlzxtmHARm
7PoCFikvnktP2xXvdqkBqxRkD3J7gO+1MLS5XxnyckYbSbsmNcB5qK3lxW32HgrD
dvDh3IRrwbjgA6vRf0XqbsAHC+DJ0mEMwWj96nnkfVBt+TGO+ZkK6tk4qBlCUy6F
i6nHCiCGlXzxruN+p4I/ahM1s9N+jWp/Nd5GgdEYA0Be9smOQUB+juPN539we7tC
QeeioAgNkzGC4Rfd1Z9vGc4O4Y/Y6cQbV8SOyq7fnveyQcXZIYzWn8sL1kqqM8zc
xER4FicOh3aRL/VkCkQ2w6ou4zeo3otY0+/jJCn0YDCT2gpgoIoY2jqfZaJirF4e
rKTEJMRzPhetP/D79CfDIih/egQjaGmDJoKkAx1lqK5Sexp9kmJ3FO1h9e9ze8p4
rSMd5jvT7PCsWmDCpkrSSkqgqWSXNUo+feed5Ozje6ZTF3UeC9G8xAVp6Ds+oDKX
/pWJlxUCXtmxBN7eTf5bxm2HSUUaRiZ6VHdGEZQvdmgSoZdBUf5A5oFf9wSFvdVV
XAqMBne/SRmcdM14VMJ52neFyg3oVBB22c0Bexacl59ywUoZcYlLX/YiKk8iISIK
1nTFrbWLX0Je5hjLQik99bks/ndVQRoNqOYJOrPNPAJ0MrlbshJetU/7aFhU2/8n
F+8KAGHEQesL+JMtIbjmIErUqq/DZDwn0dtmvJyRNWNUnm5TUa74m3Rd8CexW02N
Nu45QzKDZigESEa/fYpc6xvyPJqYvhGVho4MpnI8PXDHpSnupDmry7zKlIypa3cd
9EfFSf+XwY41kg7pYFvxQXwL8/tVXsK2JzTMqyymU9X7G9Dl0+aOnQ9ZY8xft2OL
MHvCK/Z774XovFOgrCoD+gKiWHiqC7baphuL3ZxwTAZIOO2coX1rhQEQP7ilFa/d
GfInWXi8+C6G5zyWKJ9GirkFa99TWyE49twc6C3DZOzUsfH9RLIz/+PfTWnJzKyG
ahcfhxQ8Nti3cHJHm0kPu2C4skO79m9IvTpRMcN2l2omFcar2iRXzGwIiVKD2k2V
otAOkYGnbCYW7NGdQUhkLA==
//pragma protect end_data_block
//pragma protect digest_block
NdXyTpFbAOJPQ8I5aA2VNPZYVBs=
//pragma protect end_digest_block
//pragma protect end_protected
