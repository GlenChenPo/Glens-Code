//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
uCLDlCBBfGf9aGnJRjou2aWFyahOGlXeH0f1qvslFqA7ufnLnTi2ps/RVzuTzhjl
FBlbswQT0Pa0yQEklb4nh/MxxvFqgrFO0cVA7S+06DkAQiJCMyR1pf2xlDotOFsL
IQfXcv4nhAMPyS3Q/2LJEIX3oyvP7xkI5CMjhXMaj9xrjbHXnFABuw==
//pragma protect end_key_block
//pragma protect digest_block
d6nGU7UwKgeeU7luzAKq39C5NwU=
//pragma protect end_digest_block
//pragma protect data_block
BgtyegngET488zR+17ZBS5aBMvxuY611RTYv7GuM977yxCv2bH3uebNJ0qNcSh0I
2kBliD5ERcggPj3SzjZLMB5mqPdTprMVky9L/bCAh9Wy5l2CetsS6fdZLAcZwnfz
jkJbgvqrsO6hswAIsFxK5MY+gmvCp3LdvsZSX2bUeZqVyR9so3z7W+CxOsIPxrIy
KGsPajyK3B1o58XD0p+rCfIBeibbombjhBL7WnP5vlx3OhqZA7q2qC++mqPDpyk2
7oexueglENj+Grf66tpnqu2Ti0XVHOkEWl74DuOHDLcPODME39+gYIkVhGdYvIt1
+OMgbDrDQ1GRk4MRv/35Og==
//pragma protect end_data_block
//pragma protect digest_block
OlIxO1mtatPj6T7BKWxfSp+XsMw=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7+05CCzooS6q4yyaj+zisK1+qjQQfjBNk89XimvWSE91LFvr6fFyXuAThY/MWRHj
temcWnVEL5npxzbuSgBMpZd2z764ahm8kXm1+HVO0QXfQv3PM7n0fcrDAo3b238W
prN0L0rBn+1fOe98rbfKWS+C/1sEuFJ+p3VgP5jWV4Gk16gV1ESqgw==
//pragma protect end_key_block
//pragma protect digest_block
oXBCYqE7RNYS9amHHDS42ZwLHys=
//pragma protect end_digest_block
//pragma protect data_block
w2lCk7xpjQzVbpLZlSqasZHS/NB/Q5ddgXcpH9BqhAKlOow4zdi/OR/s0mXcLu7H
eio6Pe4mkNFzzZSEU9J6FCayDI4To7aMd/5lq7w7dTrLpEMl0RkS108Swve2h53w
iPSbyRb6/tORvFVnP3iaTJyWwdAlHSlkgQ5ANLWAk8hVgZTa45hSaqwH0r8SHdQT
0UZVyZ5GcItfHn7jTCn3gxpo1Pj93/o0AxUAdMFXncXJLOk1iAP4yKqMhkyBYJXC
+w8Yf6x5NlcT0PKBXQIm7WHfdmz8KcmJVo9qEe4oAuUDUYhnNNj8O286MFsWR7/t
Ixk0gqEZ9jzuYgu9buNaqA==
//pragma protect end_data_block
//pragma protect digest_block
aSpU7szD5ToWuOTFDmo4cCNKu64=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DJR+yN2dS+hq9ulftw34Na4TjSYr7NliC3YSiJjzFIledLBjjfvtWFj0gOXWeo1m
BeBgtu+d/S5WTt+gtO3QFctgx0DNHoSBzcKq9RIYIpZSOa/1OGxW/oqGrXstNAbc
zK32bJA0fGd67OyoeWrwM84Lz4O4KWlnZXD5S/vThJQlR10NGoUKbw==
//pragma protect end_key_block
//pragma protect digest_block
lAxrc1CSwlAT0Fw3AHuzmoEYwxA=
//pragma protect end_digest_block
//pragma protect data_block
ug2RlmCW/95gYKwfoPTewdgPAid09gv7VChnUE8FJ4Uny1ANloVmPymaIxHoyyHu
z1+T8YOZkhCkOrMH4WJncm6odMkzlkT+Bd0A5gIXmgfilwBhs+HSnvDGKT/0NoQn
rBf9kMIdMGFpMIaQQjGMwSl8kshAOWdMJQiFVt86If03A/JBKeWVee8iWJW4zsMS
bYpY4aCWq1p37fy9RHRdkgmNcNQAUCvBOAdLk7f9BgZSK+q61jBfLf/8yl2rvOsJ
i1xeyBDyfXrLoZIYqGZxd/9LYEFR5USiDBqRDYtb1FlWmeyS7Xsyy/JtyjN+ylZA
SGaxbFvb/kvjaGH97cG0HvyvUuEngUCDbS3SXtKNgMEehc36wlaTWWMRLt/Q8hv5
OPreNd80fexOIVwQhZJw4hrSuuFwXibwHuDJGIXEYi/yTgwwFo+A3rerIgGi3hwD
ZX3DQpeeuoiGezQfKE0kbfI4oqAnTKJDb9vic4a/oAU4JOoEFfk7gdvW1SWq59by
wOVP0XtOTWDt5aNrupyOe8TgEnIlTxXjSybi7TWgKmyBhGS3UYX3y7MRtiJnZnwg
bpXl3lXTo6Ckodz7yvRV1wguljvs5rCALr9OCO+uxqfsMOIHlfWLDhC0jdRktGxn
+h/OIOeJz2TZp71qC3Jo7sSYKAFogQsP6WAA0pIqRG1W/naiTt7sB9yXUYUJGKvo
5iCssRnDZcL2d6fAG6z0d/pJRn5+RrRrX6BW+nQCNqhDQDMSfZ/7DEUo8olq8d2x
wWXXnIM0nxV5MRdMEjZuy+zOPBi63BWHEGlc+NC06kmdBXEAOCWuGUV7gBJPnTRa
Oe2NKUVNrcoBlvgd++aZPCnZgMAzHaIA4Qic8wrzb//GfG6CYIapyiBjG+JVGpSD
bmZEs6TykpJwk4sVOyOud6Yb4r30wOjoydN+NTSbq+XNNzbseKn7TCZ3+iA6bBW4
ehYV1poA7np9vdwpbdMDhB3OJZYOvj/tq74EJdfTRehfE/vW3pQo3FQbifZkPjOK
38n7vqOmId9FzytM3k8zT3jgHM+uVz6uJ8e1QE4d8gaI9/ijpSxVLMi5HJcNwhqz
4YX1H6cmBxNnqJ8+EUtbpkcRjQF710DFrW3clJLv7BfvWlnmBXGhdMg45h5UqI2q
aIQQa5IkeZXBWWpctrvKWUOQRyvu20UjmhENl66SJvXOvEZL9Ec+Z6/J0oU4EV/5
WK/QP1o4swG2DD3bNotzF4+6XQ/IkQwHIaXYyOHdFRLgh5o/YDjmXI8Pikqp79Ex
3T9oQwdrX0NkAH9l5TGJNNXC74Ci9fTVDTwzg6WxKASG5KiunJlFD6VG/0QvIri8
pTFqCZPf4a3d7I6g4cX4WF3SgrMTvWfP3400SqSaRA1Ie6eNxXb61p/Zokh/Z3sp
9IKHH9oFPRdAKelQ6viVI3qWI8GktPgwZJ/BX5M+XZZp67ekW/B3MlZ0BhWoZkGR
yrZrQ6pgQUT9ekn4Lj8sWpSAF9jkd4IU0zaAUlke4vzDaXnbhkhMX7eIcyE3Z0fM
Zj9BgBcZaULQRGEpbNv6X3vGg/onxBmnbn6yKhwzJpZGQb4clD6hx1CA1fqcOrZh
F64RW5sqeBejpVTblwVVdBFUPBpU0DeD97Nl22aqIkwEtG3IQPUPvTADxP9fzpK4
512DAagZ7RLRALvZiM08Ggj5jeFQeGn0kqn02bMYwtkQZRcqpa3/6m11cxevj/4T
QDskPBWpMPXnQ6pT2j7MI5hJGwoIlw+4UaeTNycY/D+LCywxrrYigEZSTUtF4IwT
fH8ZIpungjg7WxlU079O19CINc4lmK7Z0vRBGzDnyhnhl6ZKwyIb01ZdcuD9L3oE
Hnv8howJ/wzqH6CHGkHy1xK+v9pduarrdR5yzXe25QrUH1b86FrQsJ5JIfumrYc5
bJ3BllBz8cmyvWs/0WGCm7hxdsAXRUliLM9FaAtcyaNYlp5X79/qAZRCbM+8rN6W
IR5di3wc9zSOl16RtUdMen1tid5DmJkuMQJG/8YivAemG3qUdhzWY2nZDhCd6IxN
2hNvTEnjwcJQy2bopRMw0OEFAxVLqjnL/zgUezHxsLulM02Tf72bUye58CeDpW0t
EL/c3+mdeJsp0TtN9GiubSeM+d2wZWp0Ru3oG5Gka0npdBCiZRQhSDpjAICewEVQ
Eq54Ivg6weDBOZ7U+gN83U9lTF8Uux5En8xZvBs4Hvg53+B++1oCGwrEBicPnE5l
zJjRFms/s32DQd7K8zMZZ0UhrryB9rsbnqX+glA0CIufIT5PQTl3ZWVEDo+/aDiw
XhuELjvdw2P3xvc3+k8Fqi1ImSeMLjgxhBIHd9xLRfCZPWJafK2+rko01dQb5CWU
L0cXseyV/ktSaJ5IMP5Z5ZHp/RFXHTt6d/LmNU2Er9ZmuJ+PfuXFoQYGuOLee3zH
gq3GvN1HS2/s+F+sQfZpOP+m3W+eZugAKzcD93H5J5s0ZNipdgBiUNj5I2pELX7H
xQhC86pybQVGrUFISu/nWpNyXKKgGEeIFtvHfx0GluqmzrZiSdTPt6DMFtixHwKC
DBeOv/XEZQDsqVFe5oXtV64UoTjJJleynlVwTzMC3n7K4VcotBUSBIE+6mSTMPTs
8i4MeGlm54s2DCCJRcQrLRwm3xyCQaoKGvLKA9L/fP03Q2OKnyAVR5h5BTYqOPCh
1a2p8BkOTKfGw79Q7s57kM6QswgSfY6B/nqUmQ2w7YmV4ssJlO+AbS7vmjM2zWly
Y4p9Xm3Q4k2zM7sk6TWaGylJGGgFJg+uDD0KDYUFC9lMe8/BD/j29UGj73r8ltB5
0u/PfgjmkJ4Yh/G7FQ+KwUZVnh99sdNQvVXp6xjPMxLG5LSXj9nZPIVtYb+O3RyM
n4Dc6LaJoPP5IGzEwK1GFtJI3sfG8Kl8SIkxXf9TYZ3Wszk07X2IDwRMucyFqNOQ
S6FitaXW5Ab3V2mjaE/QK+AEvscVCqgOLt3DDNwH4DhVRrJ/+HzRVYjnNYhuY2DA
BrlJpLpDjjik4nodLXKb+Qp+DqyE50gkL5XNVFLlka/4F41ql79D/P4AxupVTlDL
UooIfQgVisGh1spViV9LuhaoMmoq6BagapaAN4TapP6YxG1xooDF3/1OSXaKKGum
YirFb3GjefDl+7oAYagDIWuaSEtyR33og1G9EJA1aWvgZIj4ElDp3eGKA95BkqyC
RkMxXkVOD7K+hjz747k9w39Yrihg3MlzAkPjRG/leUSB5s/JXz/Rpdi2NOr/aDB4
jYtHE2XqWi5S7mw3fDTUw2PHZvvNaWipdX4tFoxCgdr01gP6hK69UKaAC2DBL5b1
6CSfhNzt9WU/WPsHxoQ7k38of4vUB58ts2OZz/51+rub5aVgZKWsJGy4Erz74C2X
gJWgF14CMpTC4A4P8nXKFMY2uq5Cn9rEBpMr9KMdmnQmGQpKUOp3eR8aIhdOKrpQ
USeVX1wd6GIQ5jiPPOD2zq23FaadGILXH6pxgQ+R+CcagYHa9kNDyAsyGFpa5dlX
dwcCI38dl+vGwFFrtWMw32zqheGfsaGrTQCg+mXpv+IF5/l2JV5jQ+CCRqv5PI+2
OlDd7c4W3LYoL5A33dJQY5z/Fbn6yrXxEkZFPQGiw0cx9ACuwrpYwfSSXCX0O2tM
9cp2MIONV9c6sHSCoWPByAWxavGzgHLaP+lLaMp53+nAowOrROz6yXgdJ+6Rrel4
XpV1iKsWjM3f9ZjxcRYBvDMb7TD11Y7opijHniQnOZpLBwKRA37T8rW/+acvOjzG
px4jLxoCBtTkULaPM3DuJnhjtELwA0bTtP0CiqbI4dLLiJy7YFZiZm1xYS6doLVz
Isl2eT9aVv7EhAatKjgNjzxqA284bNuSjAExnnlMnLoXh0i2N9aQTH+clxdoWxgI
2XukJSckP6yV7yWa7v5aTrRuA89zaFZqX/QQxxa1fgRpTK9hmWX7qYXEWP0xxvvR
ghNYXGrtYMlp6VNUHiOTqY4Tj/yoU0y6CWQa3hBGgcTb1rp3iesqSlJculvl9KIy
2svtWPytX82wRe8RybUVbOdaeHSJWptW7J6Kt0e7z8w69hpEU9loUbmRFCMfFdYD
8Pv51QFlsGh7x+fyq+K9VaMKvAPB5n9n4zjFkE/7GzdQftty66Dzn3fhBr4UW1Fb
1qIuQ7CQzQ8TSCEqehS2otLO6GbGYX4ja14/xlmIH2IKvcwRzgzVYjph6tKC51Dz
68XDuwR2CpGvTRt1DkKVf7huex4BP4HfUnD7GtrH7xH7O2eNmYjQNTYjXGNPbz9D
1cpJwy5oJ9LakN7pfV02rhf9+3rJ4Q/EZqA/3bHv1DwiJX80FKHyC8crtcFcATGG
gildBxBSESUHXw1zl2gXxiGXofZAFhKNxwUMaNXdOlvSN8Vv+z2wkdIo7Iez3J8b
E3YMi01dc9w3Jv4IWTgJgOOUebZxA5TOf2ep9ppO/cHENaPLQiW33TpVhCCqIZ92
A/r9FLWwBpqJbO9q2Abdsg2EKMBFCgaHL5oP70LSYZLrzSbfm5ObMTTx0MWIcJBx
oX1aBNe8cxgVx2fJJInxWnUk8gUHvT1pYekzL10A8sdlCFDPX6VSOBbz+ucUfyHX
PomEtCsHcZZsBevs1RsWhFjBZY+VVrd7ZjJwEPdFbuHsPK17NjdbOt3bjmvPHSs5
YByCmVqe7z6niV0hy4EKsncORWMGbgSTlbVTwZfHrgze0MLgMK3mabrtpn+1+3FE
at6MHQ84FS28s7bJU5w1tJeGfUbCu/s9tAJi5zpC0IfemFPgQZSkv7kdhrAnl+8Y
0ILcT/3Odph1qCLTOl2ISmhQYWiJ+AlHlXJF9kCsVZKTHbyqUxM7xeCD6pdy0iHe
HQpGzLLq1DQ4YpcZpX4MEFBnpcNnJ2ZiXhmgPd8Uk5UDCul3KGTURUD+9B1DXrCY
6+stvE7IZYxoR00XlU3/rY0nPe9xNSnCHYEI7AsUgzxEpsNKUZIzWFCjxUZfTMTF
/6g1+U4yfCuPthesQFGSQ0plP0s+Ju2VkuecZd7RDS0rI0Yb7cZOLY80Xv4F7nc+
7SMzNiIRRr1afL6A9xozLE+nQ8Mqd37wHtd/d8iGR1+VJj79s/sNC922Q3FyJmZ/
RfQTfAiV0RlDwUTnmw9Z2M51mq0Jp6LQnP5FfqUzBgB/p9UPhG1FHXLkzOeMwhCf
wVaVa6utuVyzFvIAFU1IbDqlj9ybcQulGhg3OSqPGCJbffahA/g/X0tJRqsHxBzM
PPvlYT5B3pMLZMxpUnMZpRFmQGP2FdRK66ES2bOoCsrdhirihkG/AjsbzEBuPu3i
EqBL7rcSuPLu1lR+5jrB+zoKdo0OXunbAyI3HCJpVsbYnfAWPxIfnHp6JPOwW4Gt
HA4gIGxJIUCJ/CXDWalQdfqGChNw+hciPOfagObwZ4NgmLhgWjLsK8aCMg2d79XG
949ZrsxBb56MHE+192DOWhrh9GLQh53ZkPIloA/SNCkaw6dRTz6/3ZuhOotV6K+I
+GKKDu3nf1Y3tTcJCyVJh+sXxYQW5yzoZSTl5RWf8qh3/dbSx3Sh8MahGLkPEYal
CY3/f1XKVNenhr8AHTfZk0HLz5XgNHRXQzUUR4FhaHXxAhcldkD8GFhOX7p3sp/3
RaB+t9JdG0oHXlhXEk4e2YW6/umpwrd9TEMZUynMuauEIgL66vo3JsB7JiVSBsjH
mbMpYNVUPyl9jnAYhOAMigyamQmTV7qUWN5zIc1hdUgK1SGtYkXJ4P0MfmU/H3Ht
UkMqWYSjEwWjB8gBElmcQJY2tqBk/CtTfI8OFyxaq4DfAJ+vi8yA2od0pCG3Snhm
CRu0FTlg2AYjIvvYtnVOunR02H902LUA3uV7lFqvbykDqO7CwueHZCNZUb05ZQwu
MSZVTsC72+KsLkXD1xclSd+93lpK45KuY3+9cSUZlCWpdFuoRllOtosC0htDDCT3
KhLav5E389itQwAFC7pI+PgoiCTfEKqSpJw9iKeF0+xX6rv2Z7p7VEM3V/RN/A/J
6exoweSDLWpqA4r8n/QGzXsJ6qOWiro0vyBmEl2G6QM/jHzky1tPIljgVmBO6/wk
FB2o4FgZHzrzrKTYEO6LWvpiLtkLOpsv+4baGLov23LiADhtnKvNIReYtagA6vln
NOtJQgZQ9f9mpdN7CfEh1Qc28Zdrj5uM4x2BLiI+lbv2ecIZK6bo8g2oUMktXzL8
SJF62SFOuhESTN1d8VC9Kkw6T9UGF4nGLodQNSNOX0g9JHZwyq+o7K8Av3nx+2DN
XAIcCvKZM9FPC5GZNz73zd6oqHOLO6ZcDbtbpwGSQz2CL5U6bV6tF9uyWtBJq33K
lG/ShCBPOou++ovJF3apXnw1gYbyFmr2UTd9IE46msMjxPb3xuH2kCklUKKkaUFh
Zhq2Z5M6FLGFiQ+G1iMifIhAmbOrcXwecRyNu5NPMli/8g6ERcn5JvPsNOZv5g3O
SWlnZWH4CFQTFLZZw3aEkEb6Qim7iORlmlGGGgc5O35pDZDC7uDH//70a/NrFeZT
1YuEZxRYCWZUQxiZl9TA8TN3E4FzfLLSBtqr3LY6RNkHKlpXP4HCiTCpngyzLKQL
MQYJqv+Ip/qvioMX6ph5pGDspFgHyg4jIQ95CwS9DZPUTy8XXt8NAbdvdrfN+VxY
qeVokA2LdC353ZUQNQXJh6JJmJzXFpSDYw78Z/ht3MdjuWIOSeerztSGtA27W6/G
E3GcJDNt83R3n7Q/RpxqUv010NTFnb0dWAbMidz+0AbVqofgxEhlhAC1t7jnU9+s
ZGnjrvTzlUgVO6CYduoZ+fah0DUa4xt8ODO8/2l+Qc4hrRd1sUVeUTT7cZjuH3uP
ssTqQ28AKftR6BbUBs8I3GiLzKfi9DMfS/7qky/eE/lnFLCGQkAwjgEh3kys2/b4
t4m2wlw7kF5FVLUHJk3QOg2xEFhjCZ9mybvkjo4Ev8KnLGupnHBpQdIG4kauNYRR
/m1PWW/NzW62jvEzTm4zOckL4VaZoeQDHmHImZDlD2SZGY9jiU0eM1xNcmaDWRsf
0P2OCrNPm/LoSNOasIN735EWBXF5W8zIim+33S4MSb2TBgZMNN24IA1rQXdtP671
CQJgfVw6TjNUgePCAXlj0A6dR7wfENTFYP6IplBqx18nTuAcmmFoeNLDsrkyD458
V5v5nMpBzaOePp/VbzQ03vcIpwWqeJm6MWplGh+X4/ety9xjmBfdl5w3Nrl58HcE
SB/B9OMIli/aC9FU8cI6O1/oJnAWJS05xO0HzUFUMwrsFLXcB1xKuzEXDJEcc1MM
55rCzCO6YWt3YQhducMU1bh/USddoLQI4wkvLE2I4u9P1zjJUzBuZYPiiOztd/JO
T64zFto7lJ4lOyg2eAC7AcINdjSVsHBpU1TgZhIDX8TnQ587WsxrXA53Q2xuqlqD
PZnFm4poPK/eWnAnZjb5DMy5/IdbLzMXgdCqGzvOrFQPwKXxBdkNKW9IkBUlKmRe
OCuekP7oAmjioz4BVrk1245ZQOb+18OujF0Cd3J81UmuCuvR+yui7VfSS/O281Jf
qHE4MjRqaSpni1zmG2NLBeeV5PXxqbKJEOCcYOq7X8x1MjsBN+QcDq37IN1W1Bio
H/q0MuIYpA+E1ngZ49r9hNIATaREExSGB2LjDxFK079pIrxLE74C3if6ZHljfEm2
dxjCqEGghkmoyKoUTAKh3IpnmyJPWxnYcglOdUETorj+LL1bXUsHY6XDJa7+WNGe
atpO7MJ8aEWcUgp9CYZazElzkCBzxbhE8R77CAOOKHAtgAOWgwN/gdxaJcTB01fg
5/DJ+lDhV5/TfjfSEnHqGyzi1kURc7qYGsZeGeWs8CXOUp4J47W6pCa/Lks+WsdS
IeeyBLjSDlgAAf1KWoKHMorNdw/m02lldlLWL9yOqF8AlQ+Q9WWCNi1PmgM/LErd
brIj3c95O+5ZKk2OG/WtWqAFX1ysEd20ubYaBhUXylKcwO1dS1QGOrOaxgddA/qp
eylWahKuyc7lj8IPM6plSkr1NRNUGs5ttEuMNMHNpcLbUWtLxM+Xi9j2EiD9V61I
P19qG9Pjw0LES0D6Mn/XX262+RTYw7/1hawavypjZCr1vzjOAhj1iehRSVX2mI82
hrlM5/JxmAXSqWNPGiJ6Yy3RPvuTupURWobZLmpp4/wWhsi0xUazcX3k+KMhKDA/
cyS2IeGW0/A/yXl3S+fMYJGLUN9SSrGhqZtezlq8SvaDcFvNAJGA5ETrGzJYcbcJ
nTTXVw27IJ4REh1e+pL1NhDSSOn1ouCgES5rNLrbBJ7avDiDrkC0MkfaxT6ArRCn
FLihYiKroi7TUO41I6eYZvuljIdfV0sSpoG0n3GqT/RZhcCWi24dNwom4uRRxisA
bZWzDQMAztG2/GUQbvlyJ5C9YOk7eqPXtj8ClH9xfKhM8806Y+kEw86wIHTARqAI
iJPHO2hTD4Lt3K4Gsn7ugCok1Y53e80COySraOQHjCkFr0hg63ovjWfQsaR3PnFr
CysdEbkU4dwuAQBfDhDerTpq7a2LaHyAjzP8v6l7BZoHrdyCOjvrYzEfkJJsZ77B
la+rSqREnrfMJ7jOKNRJxF6n2s5HkOxJa4OOAzMJfPBCMgo2M9h8/saOoB4smZfJ
mKnu8IMahe/DrunkFkmKSHcgqrNQCsVB+MFCQvj2HPwSJMLKauWIKaWxdlPU9XPH
Shqc4AfykxPPx6gomWOOkM9KuJnUyZ1JxxYiPVwkpjkJKdF4LQ8p/cM9QA51dKim
zV0w8fivzmaZITHF6KE+tfqMgvQ4KLI4T5/pGljOVGvqkWzz9LmpdmIM6it4TI6E
jPHuKsMWVkz+8jtlNtLYIoZw+bQDc6PRWN4Kx6dPgVG65uq9DP2Yb+9plY2N8lQS
ztHpZ/7z2v6cwButr4SoGHOMWrMpbLx64PJi7zV41gDM7kUWhu9LxC4QPMqme+0s
ovybim6mjDD8ozam57wcrumwul9SERyTXFIRSPPYnzGZjpfv5h+lCJwAGJ7rSJZI
ZHKVkuQz7rj4ZW+R/Z0SLWVSk6hJdO6/gemzJm9XZamaoviLfJnbhHvYp6Q/NIyL
1iWCKgJdIs6ToIyAwN7KKYvATSeo9DyGXho1lHSNqTkm1ruvgajsTAvxdk5pD89A
HSZBa/2IOcJmNU8ZYYOMBtWCTZ3/CqHFZ7hL0F1so6yLGBm9gOCiuINOzxeIWWoz
Nf33U07ErDvXCH1j54bLm3tvkoAbegaeCFGEs2PC5jJqgMUVTHA2mrRFwENJH9NY
CkSASddlOhNMSMuOiKAJ6TlHXUMAHC3zT8z9y/iC+dNSOAhFGnCPCUd6iOQYzPM5
dWJ+Bf4+l2fJIv0bP6gSqZB8uBVScB2cq4l725zWxUroqvGxeHwYUyUl4YWKSVcv
H87iTzZwodnx0NWciOSW0kAb2zmAwfnVXKhWfvJiCfIZIXnYzbwN5IASmMO5RKp1
65q32P/kIv0XPxnRxgWB3HUCl9YoweLmfYNTLKltrJTaunHDWTkc3vqOzWJUVqGY
wxk3J+8M/9y6tKHxM/YC8mGDBCWdVc2Hx2a7+ksR83BO5Ef6RwcOPviKndxCRe7a
MfKpGCsuNvDTHHUtlv7K38rgpRp8l1kLgqjSQJJP0nIe0qW+/C/THtvwltkzheeV
idhR4zMLnGZYvJ9HqQt2rrZU5suYS4420+iw09hE0mzjgvWhoauUmNRdv2zFNWJY
fDY8DtUKaFHMnVQPp5dVzLKLlpyE3icS36cMajx6HFvsOa3XvP7sqDa59pBV/oKH
ZRpQ7WYrHUe+FR9eyW9LEOgwXHeGg2fqodSb+tPaVOPmliktejMGa0WVOSLCrXBy
OL7DTO6h3NWEu7wJap/e7qIJsUkBoYd8CbCsA/neyazSdNeZrqUrRnlEboggzFYS
x4g5irL3FZkDwfi36WXFSdFoc/DiwmrnZv6uUcAIkuUf4lFNtb8nWnvuNxEywSDO
Ua3SAtcz8jR7ZEySB+wJI7u+GEuF/83QrjpotTJUI/x3OGWh8ped0Z4LEKfECxSp
A9MJkeDXfwxxVMWxQJo9Mvklwwrbe4ek6s6iucMcLiCF5HG57Rc/pbO6qcutDIYc
ru854lqBO1FfWBAS+B4xWGLTBpXiH7T4x+ko/IG94cWryR0cDSdtRopR0ZrKfZOS
OWUS0coG+fSHmk1QuUfs1ynA8CYGXzG508WUF//8Pn0Q6sYuPkMwCSFgma3onhh2
Pztx6ZDp9lM6icgyUfzJbfHykLk6ZbmSvv5JW77lc+2nSIuMZWIoTTQjGad5BZQf
SxdNtb5s8gT0wRgmske8vDyjxjUxFsxutL/FvtjFMkQwwfEUSekAQnYSeqALL1Nl
rIrxk2MLeH2tccncp8VdEFs1Pwl2WCx5o6/+b1P1MMFrCYMGgXVgU2vEfebD38YW
5MoRNBamdFXJ/XhAXGNpaSjjPJPmRFQn8vw7a7NCTh6LY7DM6/dm/TZ6dqudpIJj
EXYfQl1KZJNXVCgosDs83fOg6BkLw/DaJe+dGjLN5dHNGFL2RaDqaOAuc56pO78y
xBIB8K2pOgO9YukLFIdW320qlSXPxEz6JT2b9wM7BLyfKMmZcGvG9yHKN1vyCnXu
JUXlnpEjzPnT3ddsZPXMigric6XheFx4SwuRB40FwNxQQpMw73x/3sjxp52OqAbE
AblSQC7yBK2z4dg5GbV7Y+PBgbvc1QUZ5t/TPAjucgQuSCm59Rz5kEIgB7z4mP4z
wzk+YPI983fTSS6www11riA0rTqw7XEeXtjW/aKmiU/oJ2ey2HZVXsJ/lL0PMV9R
5Tn1uXwKKsw3hl8q+BqNX8nLsyT3IfB/oJPptdNpwx+xYC/7eeAL1sCi+eJJzMum
bp7afmzqRqPMVwcYOfYfWBe1m/boYSw/E/txuCCkm97iyMJSNfohXSSGxMmTMEac
ztsUOmmSCaWlmI92V59omI6Obww8VG3Xz/aftD2aws42Vv+9iOzb5fNUAV5hfRIs
tzt1Lual0QRFZlS8fzf2AIzSI4qQjjzJdTAEsFLZSgPynjHJRw5+4M7MRgYN4UKp
mjHGNimtDFcnzXB8gSw+/QL5rFmq66D6eDFqBIussA9cVGCgi4ZXWj+3E2gjI5yy
eRh2sC3OXG6/RZNY1khYMdNcbjN0jNielkdWfLROSbVsrnjGd826Q97cfn3VC9E9
ioWT3HvfbunnEpeKtzNlnPlzmVetjUruLMCD4yFcqL6PhVnhP8WjpIh5lJoxv1YX
eo683kvV43or2kE4R7UxXDh8dIIlIX1g4beQJxXzRVPGLyLEVSR0zPtn3KSHV4nb
nUeXCZt7hRdVBASsIwu88g5ZKOnPARsiw6+agyUlBFGztLDP5M0gUfySdqqKHPj9
F7fiTyzbdj8euqQSC8LtpApdJPy/A/0RjjOY6uWDlvedkGM3r11qOLTxGIgGtmae
i4pK8zh6yXOY0fr6aoqC6UwSZmAfyFhf0wFcZTuRXVZTE8lmcOQGwotYIx4cUm4U
wNHRUOmPyd1/Yr+hVLxyWHSYjrGIBP7szK7s+VoRlHh4TmyKVWwoJszqtBvLLgu6
kds2EEvNc7v/im7U4dT7eIRdICZR3wL7DY9QTfB0V6blDX9v/finK3k7ATEMfdvf
DavngbuLAIrrcrUhfbkSOBVxrKNH+96rUnTO4Hj1q5TarEr/PqmmMTHIM/UG1c/A
3MbRSz5pGsv6UYJ61ZlQUURIfbXgYMSmtVDOA+oVDZDKOCiPHL45/rJsLWSaGMFO
L4y+9y4DJl4DEE0rJaN59LSlJIOKgqAB+GK3ryRsLCRGdFat0qw74cOv4IUyJf01
T6KlEV57ivO6RX5Z1hK8wHE/aZLoZJUv6pv6QX0djOS6SzRZBcuHIJltvNdTRmQE
wzEuWJGibXmoeqdZzhfUeU/Ne4mnLDyloKHXuNQj8plW4jcmBYbr9V80vheYRbac
ENaqV6QxwKrV9Mq2xRzf8k/qzI+wyrCJfxlIto2RWPV7zv1nXrhqaRhXQ9/yYqCZ
DrINFA/U4605b96X7tKniceDO1wOGZX96vyp+w+gHSoC/gKGY/SpO/KikULybEXX
kP1bo4D+qjUuwtz0pfen2/XcVhgkb9WEDdJ30uVqLtBecOwtik/4Evb9FcTI1vV/
3mH2mde5um9ZaTYzppJUjzvCl2NoP2GFKN1kgNHAIKz/BCcII/k7D1gE1qviIxCH
P8R85+G5yflTsmj31FY4ezOrxuulK5QJyTFAuVZfvqGgcxvtP+caNxlmnJ7YGAs5
xAsvaQlZC5Eyp6DJ2RThLAMMTpnO2VdPWfK3BCgu9FLBbWlw5RCw/MKpi3sNZz8u
sgUbfyQFvui+pjV+uze5YX1YegeD+L7ZuAErx7mJAzUhIWNSiDJ/XbcdGyLrFnsa
kfOSDBQgPTDeV6KnDzN2jQ/eiaU/fHAv0wofUcHtoVZ/498Y2zXb4J4E/Uioeg3m
os/m+gc+hMAoa3DbEECX1V/K+UbafrM9W+3QRWesFmX0+mJ7pK3p8s0rCKG2gjXD
pckPJ/c1YbyXZ5oM0hhUYuDb/vYGo9nJsSmslAw8HFuf13P/IOfE8lX7jWsx/Fkb
HRMxuSHph2hTsqhBUQS2FIzQOW7v5mrpx2iWkxa/OhWrLbEPXPjT6i/JlzyX4SBE
OOJsrmWLUsWi4WbyzGw/9vc71d6xmeyFhEalOiBY8ODTho5SesbhcIA4rNnoNOG4
hB89UGTr9P5pLoJN2p41QLBk/iil25DKwfpF8JNeX47yr9dX6X392EVKEe2w7d/Q
8w+GoJzfZ8CrBfhU80CzDfgCQas7WACh9btpsptA1FhGGm3jFAhW6UM0iAWXjbcz
I/XV1e5jam6Wz0KRMEx3OJg4m1h7l0xYTaP2CftaccpFdfz+bcZtr3tYb/2iRHw/
zNmtEdagxReJd8KQMNRlTC/1UcMFMW+RfJu6biAg7juTAZR3jjJB/5dnrzap2MQx
647iMYR7xKMzKZl57TmK7TgXW8zsu/g96x+ghat7D8qX+M7+N6Vbs5ft3q7uhDgk
No8UctHPUfmjmHqv0wcxoOURkVx3/fUuHhTCnUQissJz4rNrcPMUT2lrlWX2vF+S
FEa3vOXHLg2v4G5GBUqFw0qLQEvsKxSLzcLuYjvpvVF7RNMINU4Vpkv4zLPai8xN
enq63XuMN8FUmKJw3jA9DmjAVXS+2YyF4tn4LpFShAdXCqvh1QwdU8aKJBcCjg1k
hyVbfi29x9wKJkCa7fFpGCKKK3pmrRK7yd2mVdq0mKpTdVcT+nY5miGeV1a7RomL
g9h8uMCtVNlk53758aYS3ChPXA7yQ6yU00IoG4sgg7wSIf6vpMsOEVsRhxe++zzf
y2QXiK+R0lh/o9ZyExieE3QOAy9cqUJ2athgaSAkZ8X00Qqi05geNGyt/nBo9I97
F9rlG2E1ctUAGoF5s3rmOHDeJcMWT5gODjj9Hr+2JR+mkWVo3uAScfn6qdRTSrjP
SDjTPgLY5Wzcf9iX0aIuV3GUTb0ZgXwzwyIgC0/2hJabiCpNrln9H09bMNFqBfMF
Jc50oen8yTjCgCpo5ViiKTXCMe+y/lwEl79mZEb3598nIf4d1VRpVWSMjAx67YoQ
qmSNAKBPAlEvRidONuNWbws/16Qr6Ib0dDh57MVRhc8lMSrB6LOXxTT9/CCD6mb0
75U/WoP/Vcp64eokC13S8hxn2j6Iowz+fS2srr8hVBkXOIo4Cs9bxqBtk/l07s/1
IHNR9DrOmcjuBZgrb1oMh+xGV7RRWVpsS8k+6Sr1+MAJGpkiEzr5I+i3SGYZGqlf
Wb/d0F0213i5cMtK8E98Ndro1x5TzvX4d4vtmSrWN4M2VHr4oVrtEP6eZ0f51d5/
pioegCXdorUGH3s+a/klkJTHQG5+341d7ujduozcQCf+MEidjFk0zTUZg4n7Zjvc
K53Zkpj1LnYTD7tfosfW/DczldiaPQslJ+gVFqf33ZmktDm3YMAcrxiVMcGqqSME
l7suk2c7EmfksOO0bA3VCqeyVzDZDU0ZOH1iiFgnReDgbdaCyS3x0Yb212XJaXBG
mLaThZfllQc/qNx0USaUZBKPo//krJNRaGhsEw3p4++k/tQJik7d3Vfy197EkwGB
pc7Kjho0dmVe2jxcu7bCfH+yy/R0hmm80UqVbtwVhJDjJLUymVceyfu/Qf0+BpRr
WhE5RdFMATWHpeojzZQ5gq4MEo+SthBfk0U252TtpL21ffBfs83S/y59Em7RypKj
FIONTUebkLNVneENS0zY6+5ZvphrJDp2G39ZauX1JObwnQYhPXQ0RHgUMsExAqY1
T2kilQseGWWGCEAEzHiPKkpgEpTAd5zmfSrf9hyAniVWKpkGNwiWNrCcFejEJOO/
b5IRSJMoZth2pdmnKTfNjoLGtYHslo+Q6sarmSahutAFXof0rPk7L0G7Wn+AHh8L
lHXgGJc6unep9aZ2si+2YZpaCpNiI+uWLFzR8ZTnouF5sdFYOsaKTyCF0lz2Z5jq
1dffrllbFajlSpZwco6Ge8E/QvSolZlAsCEINCKSeGE9BKQI5IOJ2obiChfoeNcI
PtnODgKBo0Cy9PVvTjSJ3m0bl1PcP9wykvFc8D4JukjqkXmdzxJLkXCzDZTI0bZr
oW1fXSdlIEW6IyJM9eYV4+hCZ5PqhatGVo2e9s5Yhsh2LSaRqOC52SS/VceVgG/x
EIdmFrE7DrerVt27P3Qmfha2SkOf1zHpv945fk+vyTDfvnYAfO0fwr/zETAKgsu6
MGnbzvFtiC8Crw2o14DIe8jaCoUVWVAxqchmdqbLJYmXWdoKOOJ92m2uayF82I53
fyyCDBmVOnXuECY+vhsmJPcbIUdqtNJoCWxIvHlZngdExsS5KFaI9tNEOzD4xRfm
7gfS8BovqSEoMkEbvYcqq3Y82/2Jc0JjTx2TY8YNN6pgPHEgDsbRct0FOxssGAxH
C0mi/CoUDgB3lJbp11B8eVzpT9H0YOYKnDb76q/hYulq+kmkDCZhgPLSH/M9FQbP
zTjZLc2XgicemaxcBP+e6lwo9Ct5sk8ieYD53AGYYN78PaFQZDHWcfQ0YfSGckWA
wcFqvJ8u3FnwV3nYHxcTYXyAAGPS88bR6wE012Td657yFzWXzEt9adq+MQgbhCoE
73ZB8zUlFlgoRbusFuYH2j5dhmz0+9fgrlOw+Va+eAKCXlYSc15JOE4ji7gq130C
y9TY18Y85yGms8JFC+mYQ78TxzdUWVJbSO/646mHIx/VmRybwBEYdPyDQ5j29FMA
oz+zeE24lgIB+/YvG8lBMXwwMWN5djhyo7TCPPcGfJp0pV0THW+YFygC+TgOWYnM
W2oEwr8KkNcESX0a4Tz/+WJABgbyPBcnHzqLKFsZQsjZrc7FKrgzOPG2cc69v7X7
unZNKrg3OATQwiBmPCaVtd1MMkhF+YgmTTKdAnCKRBWdRxLPQONQP7VaxQ10AubL
u+TKBWMGgRYoXLD8gcZnQFOVKD7J48poLMCzq2+K/VS7gv7w7YZJCKnzqxuWRm5g
SiT37W9B/fIAdLMpmu9SdvKmMjgEM2kBkCmkpdU3ocISFM2X7OFZkZFZ0YRdNNm+
bfccW75tf0VPce/UsuBubeoh+YxoDZ5Kblcf6LdTya3dX018er+k7YdHUe+qC9F8
lcLO7bDyTwcg6iqQQ3WxAAAaeAq9JlOOWVYGBDbQf4NTi0geSe7MUzT5sSZeTmg/
0d2UBHmkOwL90GLt+R2XThF7Mosq5PO+HZ0A5FkaMlLyRsmbjdWi950/BJdRjYnN
5bDiq5jUS9wJaeX8DA/U3X4JDVKtea2670o0CISDppMDV84o/mrNDh4QF2mvpOny
BTHUlyzhfsoKdzruovljjZPwXIxAXuqf4fY2a5zc+NqMtRiyVFgRc/AJpreb90g/
OXpDDFgev6vU5MyzXY7+3mnZWCKREjs2HhAvO+pb1Cr6DPp50fEO9iGef4jzEYlL
MfnODVYUv2Izh6Yjf57jGZtITP5N4Y0AzrdWmmlktvYnPzelsomcoKPZDEJaQFs5
hPgOFey9baux2vVWpc2AIFcss8mRLgSTHeMtYztplMqkiWyQna5ElKFUQ7rAART3
KbCMZTeWSPnG3Ha4fkFBJyAOZffElp5EOfzAIfMKAHiujEwBuUfO/KNyHSIbFJIM
ktKDjLDgCOxgaCuoeQhkOV+KK3mxMynVidM05rWaqQhkIHDO6pdJQLR/iGAKXzr6
QtsVLR3RwlasQnw3dlayk1daxDeyuCEvku250rsWBTt2QncrMXo+h3trKbuPwvDG
VCIBFKfl51PEfDb0jiNwF3Rg2Eu+jHNmMtz9xP3hw5xPkn34eDOFZZT+jP9xJEEZ
tGBPhnXoDNLsLkbk1Wz9C2PrP/Vp1glQJVuf5cL2wNPQlVR6DfLpXVJvzHp+n8lN
hpv4PoM1I5pIshNyuaVaaps/aOhDXkYSPhsshwns3XYj4fRtUBgaNTcKXRK1/xMY
/bq3dfsfd7SYDVehl2yOcwTHTjfR7j2o6raL4hE+HU6MmWPTnKI2/FPRsByHtT98
LMJTCI871t/YJOdZV060cCtN39TBO7L/xF17AQPeSwBaRrieaeAtziS0goa0fLI6
lp6tm2008bPs0nueoOOVMm+1var/NOYg1XpoMOItUXhRfeB6W5P57pItX0d9MuGH
L/IFubaDPqCgNKtQrSIvJ5S0HTm0vlvco+M8Ug6FMa3Asc6ZcGCwmmXrxgPRXiDM
RhWZc5yy344ioxJHcCNFPxwLbMXJbVe1XNV+qHQ2GW2u3V/KsYTZza/gkQv1CMuS
bSR8d2hCiU/b0jh5SVR8upHT4Nc7qRlBfToUjRfs/SOlfhS7qLLMVpbIsLi2HvkT
msEFJB2X3UI/6DypSXPpJfy3E1fiGP1Qy7L7g5zeutjUZWISkqju01gmRI0agant
9powAcZ2EX+vQzqFV/qN9IkSHqUogytcaKrHHtLQJGIPhG9ZE3AOiafx3V2li8+k
sRVrHuxi1y9Hxc3h4wmHi+zDWmO7ILxU6614ZUkpbPJldE9U55BMq37goN9Vg0mM
ClWUaV7Nj3jltPuqjFqI8xpGyaaykoCIsTaVIJYzc+WLXDuchCQplfNUvkGcxxES
VFfmsj+/p1HQaQaAjrYkSVEglwnsCUjkPupzIUTBy1dbDY7E//Xa0H4N2XGBjy1Y
nvNymnjAUecXI9Ro9dishZQK2CEUYxRwS0/6HB9BtV7j5GsYv3YykTi8GpQiylFJ
0EFlvIWSqeci3NSzZJ9Kb9n3ILfGAM2yu/pIWeASx7pcN02zSA9+fpbXaLTCoxht
3LMu61lmROF9X0nUxDsnJ4mBu96DIMybEczm9zyL6mVQuuwNdjPWy+DJ02lWP2uC
EGXCHZaJy6u2iJXSLzpLs49hzFVOKUz2xyvmzbXrWH6Ahl5k+5fEfNhFPqmyO//E
x2FexTm5MGUyACvJoW08rrdo1kq8Mc/rSZfHMXHznt8wOVFtyVqsa13Vc//5eP2Z
qDB95JCvuAcGvKQvZa/hZwubyQX69FgUv7brgjRDqUFv+JuXxAt+aQcunt5+eE+s
M/2qAr5u74P2MKN8MJfSdgD51wGa2GtOKvD7M9c2KCQTU954LgVx/UeRy75S1Rl/
rMKhjFgEdONXm+QfLdwXQYcfP0yBVeTr3RNUEcVNRizwnRZqOt8vTJz6dG5GGEge
buob5MiPvqBCucs8iH565MKaDz6yXIwT3c/zbT0Ph2/lyCAMEMvofthAZ0SHw/04
QUXH8XbsMbM5C1Uzts3yjaEwBJPBzMocUGIy6CYqI0vUDHNDd07JvYr+t+iqssaQ
typI2ns5zOlJcmxny4a83XpI3qtKm4ZnVWmuza0ZSUnYXL21uUv+cCjibOrsQLVe
3mhUv3DJ1AsRDC7bevITPjh8shHfeVmg+ifvvL/EBmCuZpzfm2AVswAwVuEWbyOc
J3+0lgo2ghmppGxnjOjjpcITMKC1q6gcLjBF2lB0oZfGXzGb+f+AKG9wr5mQ9IbA
gKz6GIGkleGGYktNz5JiwXtuKfwJ43DL7kOqp8+oL3hfgBAyv51tnWmzaYQWXcjf
v6ewCzn23wgSTWpzYoCmsuU1VugAgwydiu+83ieTLgSRC3BLRq1hj/eHqP6houxu
Gu5fZbzWIlEy8HHtP4f+RmUis0OY3DDiZDRJziGOPg5+kMedL6xG2+RwIq/pKGGI
eiRJ0Pz5pF0wU3unDD5zm4pAbwN0ItuF1FdZ1npn3c1ex7KBf19eJBLmYg0ZyNp2
gWuuxQUoZXhm9TcrBExM+osDDtsgSLS/kIKEcx1gBcBsHhpW0kQwiIn6Cbb5Ysr9
Y+DYNUFS++5I4bioGoqoFuSQQB5wSaLz5sm6ZJzWN3mSkw/UqpQIeMVynMI4gJFT
7bb5WFx5F+QhWMA7uzWtmGuHONqizrEtJqPpaHHUXM79K2/ZMrxfG0nX3tNTvb2p
pWPsL4SYNNWt2BQI0b9v0z+JOw1AUM8QdgHuD3aOWyfrnr28Lh4pkuzgwH0NzskM
tVqT+U+yYwWIXffDjvpToEHY+5q3A5d7h+FigQxTYNlw5o3Onv0+8NdAxF+oInaC
PU4bokdVNKEsJFeD84yxPVC6LJbDrRv3AGJMslS2pXmj+ZYHAv1EEVaoMIe9f5tC
OiH5hexcsqkpMdz6T5YtHcoL3z/DM6aa186RQ1M7bN4MIMRipctMtUUQMWvCZEyp
Y506khzKcFav6TlDo5IArLYFMZITSte/A/dewa7CN7B0b0eLh6vzaFWwuhNmaO7T
8P4anL/a+a3nB9GrBkABZRPHRk2PlGPwC12mn7wO64Wn+Q7vbqz7tV9XueSoXslV
FrejXTWFQnSnqrDNHiruNEEg7eLrP2ZaNQcH1E5v1HKRfeH7Pfd62hjLF0mzIo58
6qIhXcxnycgiopPjc8Et42a5mhWe8aIHbihnYgzjT24I0+JU7EEjksLa2uGX3uvs
lLfqmJygX1WcPSltJt8rwN/qqRUHFttrfLUP42JLgVV6qhsuF8caA9H64uBWMHn+
Ld+uRvHkPBts9aQPqf86H86ypfENQNPym3lId3AUZHZ2jl54fxv5Hdvog1G7Ttiw
gC4/o2EORv3sCQhiD9O7OnnFq8sryvVgMJToGYHRkhbU3G01N1O73ofhBHebvqbH
63pTy7SVslEFfAIAo/3K8RNE2IuUaM+TjP1m9SXYaa6K0cTRIAB4djX3ashPaB+a
3OGAW2vckWPcOUIAWr7FwY1v+DoCsmI+Q5/ixxJMZzsAwRYgfDnD7iJ3s7z5AiSC
AFFD+rIR8wctdYqj4l0VgGtu1YEg2QmExvxKMlTYU6InprivQ7kidPDZsS/Eyc9v
jTJpFrPR6b0Hdzo3tlYYcS3bUmys6KlTwwTivawxb6Sqk60trR9oUMDE+EGUiFN7
24sMsLSAiA5zLioRHOlS7rpXQDD1xY4yiaDCKfsilUhgwwQUAFHXY5SpXIfWFp6F
jpFZMJk0wACLets+royIgkyv/5P+G0EGW8q05DqrnaH/AnA1CRNZxXagcmE0HhKf
RjCFaSpB5YfRzJQ4hgXhfauEEw50u9ZkCkEJMG6JyJaVUKnGi7uMN/gQIY/PUpN7
YvRbXrwS4/r94KLZip7kdLGC3LUbdxjtZam3Gz6GXJ2EbCeax7Go3yiWRV4WryOk
rsFmYZTV18J3jRGt4+enpGTWLzETpyLmlux0BkI44GbNywz2Ywaa1wSJtBjyQYHR
noml+9bVtn1f/shNfeGBRAbp5vXtxOSaCezuQXfOln5Wm0r0BjMUNaj8HYVSyZJV
HFNqadaUIzUxGAnOVr/kEoPocS1nMyHnFe8oe2Xd5ZQvbAGEmsE+bO/Utse7YGdH
+wFSzJX+hc7uOy/gR39OePYGWRyUJvzh0dL8Rv+T/+c14wXammFglTqpsxDHSb9U
CPvRvA7Xv/P0quuFLuN5qakGZvaqpyO9Qhh4bdFQT0QeGCCvbX9/Mnh2x/KPKj9j
zy/xxSmldUEaM4/UgZrLbu/+gjnyJjiAU4WxAjesCXQradDVNJZcDr3y0ZZDcyvk
rjIBfM438FfMSALgwQMXkt6is3CVry4kGaw+Uus3UWwJjtaN5r9PyYWmMRXsBxas
/jAY+BPUFQh5Q0/eBzU/93tjMloP5Ugu5rlYX8baXZSBcyRFoP1bH0qzY6WeD+m4
jq/WaRS6tq4iSmVSTroFXz8gEE6t7NU4TM/TeQJ6DbrgrEw/3ChiRILqYr08HmHI
n2CNbCkwL5zgVWNBcVrC2FyoZ1m5/kWuEndDngXTww3zWj2ekEm3+fTzllR96jSK
k4kA09eb/LMcRZnG4qf81Rg9QH8m/cvaQtS6NsLASEdLNUk3iQ//56jp2W1b0fl9
+qmhHNc6sXaaVjf4ifqUlm8Jx+EiDjZVQgYG1n/N2qjLo19uH99+CW3KqSWTce3/
x0PwuvmyBplD5aKZ2/bB4Q3QhGxDr/FU2iEtot3ayuE4NMGkcgGV6+sdoNXDenO7
KDHZrXvxGHfAk3yuZ9+kHWzEkkbIs/X2PHNTDme9ty2F1LUPtOKVT39Xv/xu18cj
ERvzj0STJoFMn2ni9I4QxKjLsHZ9Ru4VEzo2/OcbC3NtgBy/DKqSxEVsVUt0pg+u
jbfHjZx3VK+yF+Yj7+WoJ7BW5WKgtfSgxZi07B5ovTK+W/0rm9sJ36zZanw6Ohfu
Ac/SE/uVDduYU5BYddCcvR+s3ydnCLdujgNGUIBwamzq9E/ZC4WeDBzeJ1OY21+7
gjMGxb2i53WsaE2Ae6Sj7WRjKQmaFQTBHCVQA8TmmEn/D+6vTPuDKr7adrJeK/Qt
6FEYGQMv1bCe51A12TrB4sc9GZxTs3BHwBXNXGdtjxQNzukHSC6Si/hfWNEw6hK3
TjsE7clfAxwABQCR4lf1FwhZZRsdT7vC+vo+bKRtQRJwr6gSSJHr4qp+1He3a+SQ
vkBKgEIxfrp7Zgz0w9GEqQqzLjMUQFMsADa5Guhh8JwdlsjNQPIzbyD1o5X5yCQk
PK/eKqOA4g9HV27yFc0TclXP+IKqQWfZ6YefhWQ5aXsv+b0FZDNNUI7W+6LY+zVf
Huuij7dOTnUkIFs5zHSmdI3mQUOpva3S/nIdyx7KWqZFolEXHCrmtiyzbt3nlaS4
NWDFrWlgK1ZLHbXP3d9pGhV6tyI8I5LD0GiKkReuCeDURjXLowBLdgPOOx28Ct75
Fc6HcCVeW4STI5s/kmNPQjrbl5wRHaD1UQ1CAMzhppscvVJOlwRYzBEV93DBfVMu
LjbMvzv2+BPPJDAXD3WPGSZeHDWWsPz7W5tLNWp4UbsrwNNRxwY7faqHTvUXCtgr
SRbFl/xxZyBxtL+vvSxIrMnV5N6kGiFxZ5f4WIHsKSoyU7WkPFsFKEhnNbQZYrDS
fx+UpJDTk7e50fG5u12kH+YcoTLNgnXwUFwMbi7hgQAMCD8CfMh/jWhhWGTjXMWe
mlv8yOsWavMrnKE9qcFtc0N07Lm2QLgrL3/5EeyqBZ3R+czeUZFHpsPbIAKVbxsc
QQjD6yk32XkGVZSQgMi/ITMHSYMgRfQFW1vPzmOJ85Kx92PW46FbC95iJb7r/8Lx
nNvWGXrk2YHKFykfZV5DsnqwbkReg90ODE6p1y72VdVvywPLnSmxaMIHMOHwdVoj
64yXOSVt+ccn4lzaXaBnRrZ/eTj77fhItv4bidUYXA1DGx/xiAU6wxdicLhAdEcO
u78QK6/Lg77fQdxr9TZYIXR2ZtWM/IEQHEF4bQ0IrF4N8UBJ54egm7D7d5YhK9LY
Z5cw8SbZrYdSAXMO1LmGPk/96D9Syr2ROtKPogIDX6g6T6FIyJ7FfupuoDoBnM4u
W0e2faEAZodpi0WktGSYcYPYi5APfiJwpciRPFhcRW95ReFhzNekjvcvzujXYv0w
90x2YodEtIGIpxVsXwdqlV7z4XmzsK9hBVXExpSvIuMMqOECGLfaVYn3P0cFH9Dw
jSyoGCp4+dqws5ks3z5rrZTgFIOnIWAt/UC0Mt+0Dbi1r+Q6z0ljfpjWS/GppNC4
H/LCSDqs+BU8361TsbxAYPohfYLIgR/y+DMhP2fajuk3fX5pfp72hYbRXRdAh0se
PjgU0OkAdPlulGr0mOcAS6Yql2wtCwxhN1WREUBDGAUIlzHFnldPK6deYzMmLQxE
evq1hVe0Kb7ryWSjadcsxA1G4umd/NGyjnaHQhhgy74lQB0UsBIdcHvP+AfC48Sd
X9Zx4r2r2a28etz+by6TsWxsQtCv5wcuQ8p/RqMPGUKTFFdZAWi4eAl4o71gM87V
j82An8F6uBVH2iVvpLosJ3jASGE4iWAxSSLd9Q1Z/7eqsB1+g2xr8B0LcJ2r03Qu
SXbV+eobDkU4aRjTeY62q5JmSjQecZoXwMQlua5CDfzg+nKIaoNj1s5zy1FdzTMI
+GqE8eEV0BkrsGl3uTqVGireZ1wmXf/toKT+d6b1D+zs9g39pIT4xqMGR/YAKYoz
/MYpc2WhMdeBebdKRudRJGHPNhi6q3vSKrB52MQXhEPnbb6uxQVdi0Wf3jgzkeFL
ZKfGBkj+SuZ2yObCzncA/gFFWhnVrYEJkEdwYOXB/DEkCURHFIMvBvpAtvwEWx1O
lP84VFtjml1BjNme5yydOg4/HokjHQJa4fXhAe22IkOBSBkEPZBffxHDtabmm0Cg
drLfHrJZrRaj2In5Kj+h/RSMIZLoE+v19/O55IDJ31P381w2f7PtvvGghOL0YInw
yEeJLfn/qoc7q/nkUVwikEY2Tn+pRoKVWDZIMtQKiXLeWY5FCqTILXJeIc1o/dIf
vFBzXvunp4XiInDZMzxZXZQ7gZa7Zggkggv1sJjfnxL+vlUN6yLHsAc4N6PmfaPI
LFvIYPZl2MurrDZowzkxdKhhj5nDzfAAr5yqzrJQYaIQwDXPm8wVX4DucbbSDchp
le0OXSQEcAocjzPKKsje7/5tEnMhSVqllbmbRim44efr0DyeV1j/HM//SsKbgO9E
xrxMEOdA/DTQZtnyyFGZjl2J72gHutjxuRNyiIP71dVXbmkOcT8AeVRsTgmTACfV
elooqj26kLAwvC/LYmf1Ol2mJicahdh0pi0oBkVkoD9vigUwTKpNRL8T0X/sr499
BbIEtpX7NtVQ8TgsgNDxEYqxoPdMpvFdDnWVswHyl6JBumZZ/Up2GZrFNifkZByu
gxX/kfUX5RcdmbyFUh3ayt8F4jamFR7/cr0evLW85p8v0dzY+B/QfLaaPevua88D
83ymFqUopqiiF9NEzqmegspxtJ1QMG/GonuRvz+s4u9kId91w+iWRzdW4pmu4MCa
6QjgxuhnWqVSDTdNUkWoA4w/dYDlzB+CFIhRwyX9lEQP9PPPVdkv0nJJS5SuQY72
GaXX0aPCvXEzCEEE1XWzSacvOrRC3n0IvSOhwXaNCzX86Sz/G3t8fJ7KDF+C7Jhs
klqWPti0lVeK1hp8cm/BIDSgtzpZtV2kINt7wJ0Uaj5HFVHVll92a8q+5tJ+CXPr
tLFWN32ps5vgqcCAZnP5cA0YXh5288vFIIPt0yR+VFQrpNNpq7EGGA5TtuZjekEK
nzxrvtoDcOkrqRLPSmG7KZEPBMr2trkJImPArEsX/eQ5e1U9IIpQcNr2z2IQmf+p
AnSbnDaQ9EmxK+6WMbvEDkni0rRmQBE8D9NQ9X5Sc1HOliXqQzEMmDMG8DRMEu57
DH2Y2SqjStVJBdbw3Gz3HD2dBADIe6qPy4bBis7T/VDQp9CqrO6exXD5Z+kW6FtL
ToZnWEMwlZqVC0YJteKpvsuEI0YDl1CQWRZ5EY5H/EWVVmCuL5WAKNacbceY0WpT
QwetpkdtWCjMbRvpFs/BJEyAm+cB1A3Us2VJU1Q6Lqaw01RGtcre8FzgCnzxjEu0
1vnPlOI5mTU3HciTyL/tDix+nU+H8UnhxXJqH1sl7bZJ+6OirYlwjucZ41I2301S
5nrSbqyAXnNVT9MgQlzXowlxMNWtGMaISNROrYxfSekGE+jXpJhog5g5x79pnsHh
kuALS9ODPzrxcDTUu0DNb4PjyMRLQ9Xy/iqVSKHOD+sELeHSGKfLtgKZgd6vL29P
vq9MaybOwQWGX8+tEXDYD36iMYtrrBlhCUWFhYo+6JS4VbB/4ahtut4PlmwZLoVl
rXzbwD3zLW7SiL4nxxtaH3yiR2Pj95yy0YfLaQXY9Z8zDfIbpgCpACBmeevUJzJP
yu3h+HEnGQ5LQIH50IKEF0GTImV2R0Fhng2Pwiwjj9ZDlFA78SCGaBw41/O1wo6W
TaGv9NFajNpBmvuln5GZQvhCkwCfxFOY0NO1JSlgCy3SaGkHSyPNMuJ5sNpo7XFN
fg7QXgbOEAIxl0YnqK8dULFmit23J+Rk8WYenRT8WJfeVjPtqq9Z7xngL//8YnAP
905lLm6C9cUffG4JkGbQK6e4vVj+aGZKe7xVxvtFQJiXs2wgHszOyN9W9lpcioii
rbMP7dcWGi2IWBZck/vXvncPlm9zZSFFrhXzbjFnHuWHdYod44orWYF9DVCQSEyT
yrHll/+RSzlmR+eIZ2+cYupdRxveb2WoDgmn91l+LD1JVa2QZ9+ye36ZiEysufIk
G7jsvl35dpZAL917Dk0DZP7r3VoB5IThbW2UXouIvtTo5q0jM9lgKaLrVAi6ozL7
xlMsJeti5KmS0OBW/2tTmYSt9sbkK1ZTieQNnfRE/kXEZp5uSmay0Tagfcv5okre
KUv+FADdQoKj1G2Uau15hKcuiZf1HPQS1hrs2Vad1ejQ8pdAaa1pDkjpPyGffRDa
FgBUa6qbCFyaPPHJcmByC0mdMcB7ORq9hrBww88ejhqwPZNv9etC6dsg1xDh+0Rg
auGDkCx9ziIW5ygHpaLIOmW4H1Rt4LmW+7W0BS9us4EK63iGfkqOD2fyBjQ6kX7h
L064rOqV7El5pMfWpCtsdPRXN55NKm5AY7k8OTTxPNGlr9NR9fU6Qd20T0OxvtH9
Ic4iA3WXw1a+9cXGdWUyOdgyUl/3OKOKnhodzTQuWcmenUqiGM05vmcqj64zgtxG
ebaeJkTGdkKzHunAem28LaW76yggaA6CyFTAzmwfIVQk2ItfWmYf3yCPuXj9w7vi
PozvUepA7Eb6qhw+qV6VLKM3txhbrzQG7Nq0BKGs7xIQuNNQz3DjUwyFeoDdPc5C
oA9g/uCVjYYPYPkCDQ++bZrTlZOhodM7nNMFrn2O0HSH5Jg06sqsUaNN2Dbgpmnr
kX75vZUeRpRXaRUPIEU8Mw8ydMtw1hZ/hDSQm/eJT2Bj4nNCOFVQ0fhgRL645R3U
4swhR5r9EXHIOgDE05E1iGYJWuFOWl3Nz/zTKn0YpWc7mNGmEGzxCDFEx4dmSmxj
YNowkfhLrRRFeCf4vsCzE7ZjQ9ZPe4ODIiki+SMt/XZWXH4nGH2t7Ts4/zhqgvZZ
lbkurdeJt01A7E4uElvqZUyb5tB3Jte4twoKGHLnH/F0UME0W/Zthp5QcRsvEjR9
GV8QV0tsB0ek5Il0MEWLbkq+F4Naq4zzbUXUcBmgtmBEQbo0974YesRVjrz3umKT
E1pegK0BKMgIrKCVU7E95NZxK5mSQ3k+6AHA+i46QFEsB0kAB8Nw2Da6AS+hHlQz
GZVv2cAn5CxS6HhzljEnY7Yfr1dXcAopclbtvdJLpYxMThiBhEC7QPbo1rRKB7kt
1V3n6BSyEgJbMFap11in7RZwKCOJJH7NFXlNidx+tcNC5RzhTudg7iCWlHUsT5dF
kDeAakWgypoqiv3w5A5zluseXSR+qku6EUYKAll7TdWmVVPpskJOKEEhnojkkLqU
5xtJY4KzQCYmtNwtG0oSf3MnXfEJ+4NBd3k7EP6DpXiOWdO8A3BPkW4zq7Yy4+wI
Zp/eVIt6zpAJD7ZesjZ8UouEKZB3oFTamRh5n9gqHuK9xEpdlh19bIR43Fsj+x1w
Vbc3XAJ9n7pDpaZTgvX58dCRvWpKnH8Zk4dT+tbjLh5Ap8TAAwRfZTLwkzEEPyPM
bVuAd4NcRL0hKOuHDvty1PnHLIXv2ANTanh+YVqGkmhBmcZZ+uA8vf/e+7f1y2Ev
nm3rdXMrTYsxsHzlVwBp7kHQ7M3nBE1sXXyL+otNjCY7wBwIGdhtCfML64i0OCAA
8ET3xBjb+xQEXIT3qlxscNC3z2Wv/XCJbnoM8YmNt13FG0N6RDoLgAEH2lHFCNnZ
L/ehAQCeAnhIu5dVnvMF4mkOJw7pwEKDjDKPuh/xPpI2O3mO3RkGjiZRYX8MbWrD
LQFR7C+hGh93K7s3nHmZyzlyIVVMcNL9x9uCYgzEPNeZsl0bh5wqie5vPUT2rZgO
FGb7rGXc7USfDvDKyw4QNsVhlntOZihm064cUSeD4JgR+WdcDKI6XVlgCLJJB8dM
+cNwFi68p+15t3V4AvqIFF3Z4nVaDNyHqT5qDuKutuyKL/JPzfa5gFZFP+4Z3aHL
Z9302uP9P5zG538J+piDhoUuW5kvnBgFSipcdSx9u6LgSluxgYzdIbrAq5pUB390
V1Re6F+LHmwdCWzugMXiLFjtM8I1BZMNpZ1xr3s2BSeGDk9QZT/scG+9xUvAKuat
m1XQVUtbup1PCDPy8nphODIydHMPTiFKxyFKvYyKpHhfe7eJWBe0rApF4umLMRJN
YQiIjkbkVyztx7YYTWoUwod7RT/GJFLxB8fOcgYqTE4Nk7oOSa5doWBS901fnjIf
LSzX6JJ2qrY93RBasoxLZOUyYAbuF7DEkqpJbQPLxTnfNlZj8dL3sQOBIVLZ1wzK
7zfoQ+rR3ooT4oJTNqnCUfK3FAaUaEm6rST4471mZ2iKEWzZ2bF+8iFC2OwOf3DI
9Q4Z4uRscIHqCBO9rwp+Rh+PHNVz9lBfQBEH95GLb6Cy37pEk5/5MgpPjP/NaoyD
Fden35V0KVpZmrFO/f5o4n/AeF4I74MwA2hkwpFBKNF//k/g7U8M3FyJr99Ksuim
r2wz1PDZCmMWvFf2sQv+wLMZabx6l9grLb2pRGmdCHGLUXYanJ2DF8rsB8CM9ooD
rry7eWeBoQCcDYc9vfd5L1jGc6snR5Z8zrcIg8id9EdZMMdCyt5I8Vzk8agHrvqZ
sEkggMl0+VK0dEOtBNuf1/7zn/+D5+ZB/cmDQ1GgYwKK6kc2WyDlPH6SMXK4Y7d8
E/0U4salppLF9QnwLgXpMbAs9lCQz1wGLFDeDmLKtjtxDJ8OVTHHFwJvmWJkAC1T
qxbEHH+o8Az/Lrqg2oJcpZIYcKuGj94M2jLxQfK1NAi1+2QrGq8+ARL8ppTul6xC
z69IfyhMmWr23wf4KHRW+8DIgnWPh1LN+WrX+tMiolBP14tefy6hfmDUmDd570Db
QVfcNJ7/9KiPVHTbdORottLWrIrWZRVnD5OSwxwAsMwXMpFvjlJUbeuRG6AkPNZT
tKiVn5k7B1LXf/RIrplWHG4By6ep3a3WWM1g7C1TMRHp4VhVPjgRb3as7UVMUFtp
lsTmXxsa5COCo877gKwqPb/JAaJhDT+b86bT7pfwtD1FpkRrwB+697HAbZUfJDxG
8d8by61aBuHNkWJPYPWUxjuO6ICIAa0b0UaPHN62EzFHyW0DTR5yyGQsACiSrfle
TFFFrFiX7H2d2YAk2VD45r7wfJLscLIUDgZ3jrckZt5LvTJmvn+bLMqkZEJ3cZWN
DsdGty/DP91CFjrAC0osmrg26zM1/5W9aiaXvUCjp6DTZhHCP8zivRpGn2P/EhO2
+0tpqWYfvE3FbBUdO1YhK66f72aIwIj3cev6r6Zfd+u8NRWNgWTS3bh3UwUXLgIG
Ghwt3GDztScPGXj/T6Y1I0WNbakOHv882cBr6CYRC1u423YuWCuB4JmB6Q4HX+Zi
6dF5/IXlDWC7oaLemQng61uB74q1CpBomyNhtLtfY5sKF1M2q1w9dSsfg/42PDMb
+VxSVuEXzESFVshkKe1i/UB5RIClsC2WD0tbkucOlCX786snEZNSOG3Nalv6tkBK
Em43vwG1Tzz9msXLaGUFMzNjWYpT6L0tG+y2IPB2c6LazAUYsxUi78wfxaVeqips
3F/mLAC3V7ljJ0CDXtj/qsL2JyeUic0oiHEyd4oMChFcrxVfBCMV9Kd+3lr1pcB+
YBkBN3M0Z+l2MOZz9hdNiSOxqUNeESlluVSYPGsTjdWXSBIyBeJQmwNNtuO00U4Y
Eyik8tVYsTzRY2vA8leR4ceAUxHdEZ38sZ38u0PzHugtZWz42W/0rVnS+1uVbBuH
hEvKv1OBO2J+v5MoOdKoIwjnCRJJgUOMJY8Ik+kD2gaaXJ2h4BzmMZ4YiGeVYqy6
gg0AMBSvd2G4L0MezgeUAbKaD///7w3fcMePwKuzf/GaNqYlx2y2zSBvCr0GfnaO
WvjVc1iZvA0Sx9s/ReUk56RZiSp/HnAHM+RkLDAY/KdaTvzU3XQsLFK1zOcc9UNf
4vuTU698ph7g/XleqNnjYnOwbG4aVmgKYmMkTcBvuUORRv/idTbmKmApZLayqc0q
+0HtKLR0jbQGv1rgF4LYGwtuuYFNJgHFjwlkbD9cOQRoCETFEHkrzSR2GVPq6e5N
Aq/8QlujwYFyEGcH2Xxs6qgJ8JSwGUMxWwYL0NgJgCY1as6PSjvQtKHp3EaNYj7d
0q0xsSmhKk6oyIi586VaL8aAA7eOyBuUQok5Jfft9vhjOHgLiatC9GxN4wODEWhJ
2zlUscl3Z/4dKSX2wsEjRAVtLUcZDXPTHq/VhHlZO068p2EQ4w7w3akUZZ7bRyOK
5k3qvWyL1oohOEF8OJ4PsWTS2/vkk+JiBY1od1XHNvI0rEc3tgeZXNp+n0bFZj2J
uLdC/T4s61Ctiy7nfFfwBaAU1kYA1hPnTwG4Jzr3hsIqFJmYRDF+x0YDiUp8Rmed
/3v9U2hSxuy94u76TRfn2CCpTel638FJwibSxd+iPjSe6JZSN696IKFHhHZkBy1I
+oDlXfjcvYzJ4D7AJt4CPibgwyOlkbRzNoUoHNFguAy2LVvvFS+5y14wcFOwbEiN
Jn/XI1wSG8dH+WgtnrexCUTNqJdvFGypkt/LmNl2dxGYxR1iObe1+0k97yfYMVK6
XlS5lsdTmqMenHkqtuBOVOVyujcuQNomlxQ7To1opPZ3vWK7bB1bDwtZ8CyJJz7j
kxivSFEYgTYPHcsnmm7FTXY1s3g6Sttx9jUxtCSEGOA+j+6eAzG2IKdp5G2NgcZX
FKkl3qQ5xST2QJXRjLnLhU+RCs7YOdDEH9b4Bb/n+GLGd85YYtb6DbWhoTur58jy
AEI/w/RvVB1vs8UG2ifXE5SiTlbU2pYKg+a3bBtyfTOdG08qky6otwv8N0e/DCwF
DVzWqK14vIxrPJegryFBx5lBV/03iudIFF5RPP/LPy4z0/hZyY4T/wYhv6eUH+6o
eG+Q9of+r3W+kovpiWTFqaigSKzWZm4YRMdK/C3bWCgJ/T+iYjiPG3XGDwrbldwu
WqqpnKaLAyMsVOErYa/okWsaU4xFCjxCEqLqW0tvMifqC4oIDsBLX0Zf82Q9gel+
gWn8XB8h8IL7JVTFILQJiOmuIR5c4N5QqXJFjJ6irmLm+LbcdwvZrdin/F3naIEC
BECAcEKPGNgDOmIOGrG+HFR7UeCK1J2ioq3nxNv6KIVdmH9ZjL91+xw1jTwzVr9W
13MhTAGzc8HdVXXzyojrLLHLECQTiL5kOW9bfxgqJFSI+W8+JR0AGAE9ejjot4Lz
mq6pDOHkd1g00cZQprHv1ma16naVXGGllvzoa8YShqeFa0vqWd9fd5yQdEi1zKVo
7+SZwReqLBAsHh3Ug1eqoJ0b9B0j1/WlfVv1fbcBq+R7jSGLyHKfDEcVoWTUxFck
cVaAfZAkcSsh6fEE7BlFuXI5ulIrB1Y0ltgxUrUP40OCJi3AesilIT18Z6gbV9HU
htfA8mcnnP3Rsi3H7ROt6VpJLZYlYr2c2IKP+02MrVmQvtizqqT6ORC3MsvzjArR
BbwcJq06AEa7yQBnDCuxHPEXm1EnEIyksCrpv8gI4NW+y2hF3zePIQlduvPIFmKD
0NzOrllNV9VhbYY6DJAFu8Pmv2JBkGPV1hKwvnTv0R0O/Mr9CJIAi++1proFLBLj
n/hE2iAiI5t1va5+ccjzNyz4vXj4fV/scZifZFR9cwUSxVIaE2K0EcJIEJS+0l7A
LEiwqHF1LN9siL/a87LMJl+ae4fgTtAFUCOLoSEfP6OdrNgErxIUZ3b1NnuttkqO
bUGl4/BJAGDXkzlOe0FZCutRTVxrRMdkje97ulUrCqenHX7CB8WypQfKdnVIfsvS
9XCVMpsr0EURTGAkAH6cYOdwkQBcdEYppxT0DA28mBfBFxUOXeL37qoI1OG0GFwr
whqvMN0kiqiM4iVsqLJHiO+2Ty1lMMb/58isPyUEF6f0OAm61t6Vq8KpNIWARhMU
sQQ/01MUy7SMoagb9AI7+p4RNaYuD4KXPUopNItp67NtQkg3CWfBhXMPJ5FqIhcg
3ylKOtQi90NggqX8bYL8D2L8p6FhyJ4QT04wQhQUr30tfyl3jdlkKpAlbMVBIQMf
K29kJ5aaE2vdI2KP4oRO20btfA/qsrORJjfCCbFklhSAXcxl6J57edUHeNgCu7zB
28Q7/vnuXc0koPsncqVoO5t6QwY4Y8Eb+LdZ+RueofptLYI7IRioOp4WQyS93Mx1
S6h3r1tjBJboxvdBmFRc4OcjmTkeq/6O+WarnUFFI/JusIiLC9kBIhcc2I0Jhx3z
I7azmiTpLfsGLSkMwi0FIB1WZzG6Ocutsl+H1a1y3HFjlamkUzEXCs0kzTyszMbU
6/ikDlnFNfR6hJ2vZ9WV9cECWt0HzzOLVOt2otvYQD7SqS+av4JUqVf+9HRczfnc
dWX+djkHJjryVwSmzwvjfz10jdXtqAhWVpyisrZmRS9ddEM3kOMX0LpTVr9QiT/b
57+WDn+8aC4HQ4gjI0hxAtppqMhCFQJ9dCgYHZpworSGRCDHnE17mMfUjJsZJ82E
RVj+hRI41ZvRnkRQEscPwoVEwljlY/7k7Gf7a4e59qw71sHb8aI3xSS7NIG3AyFj
NHG3wMJscj6sejFfWqlAdwA1s/p+7kd1ZSgcbDxyWXYynESyq3cbFghWR17MS9vI
G7px60sUY0YM/tc8Soq9wpiRRA9CfMsPK5tAhyGO+434Md+hQvHT3mUT/I0pT4CI
jcPa/yazC1N88msXFmi1Xr/NDBbZ2s5Z1Pa34D2e3ov9jdlYdxLCcQBYpHXd4UDt
KOttjJPs3eyiVTT/5huE1eWTd4hFK+DWeK1inUmg9UZw8QIwhq7pqEpzZMoHJhMP
q9WN+GcaKtn6ZsOn7q0QrtWsLHp2vtbO8B/N4Umn4psNE1P3V9mt1raigEZQhH5u
XUwNHX521uQazzkvNROs7LV/HGmYipP03/w983malYSA25l9IOLZCKxjzwUdFB52
2XH66m51extJkIrwSXWoIbCkTQ27ADNDjoTBiTQQKjZ1bxHJjYI4kpu6jSR+DSyN
cKRNOtikSvub2qTQ0fYR7EojmMUl0qAKezqbgVUiSMjCLzlI5sPRfAkLwglt89LC
/vaRBWEldQT9OpS06My0EhksB8M6C4wh0Tx9/bbkQxw2DarbJPcX7Wrd+Rr11DSr
FUwdCxkmkMnJnwiqJm9NPtr2xcCuBhVpuPcdHMc2oa86M7NrrrrnUXobOj3hf5FL
hD3fUaso9Bmg4v5sCqN8DGPcpUfcnME52paLgI8bKuXYYo6o91BRBkDIMcGpV5Fe
MsHOwGhtSeG9vDMncZzkOTNi2KLq1E4gVc28zJfLd3bGIsVcHLsgk5+ggVb8k5n9
6sC2r5Aslu9IsT13DOp1UuD8j2y3kyRdDoy6JbY9LDVYjFJBFTe8F6EcARXqEelp
U179gpIbthQM8mRA3X6qSWdPW/WH9opOkvw+uLVEACfyFZXrsoNdvqI2vgEyaHkX
XUaxfhh+VdCZbL1V53pOLlyBY/wm/IRul41PICtK7W26VoE1BftyHRH0aVNt41K6
uStVhNlGd7CBcgX1jmCoAbTi8F+SeG9TVTRKgTt2TThUkWKP6Myn3NDOw6PKbQra
Y5G+GTpAPbfvCCRZTMEWn+EgyT1sw7Tg6IWJIFHdPZg1b5kXLGXqaMaivOROLl8H
fuXLMxWvif+k9nw2nBwnsS/Ibc45W/UFWFNk/GzJRiuvK+vnfvOzY+wcebdsBiov
GtfWu5L5VfnJsnnErfZXCQqgX21iUPoGr0LPa7mF3cz1GnG1v+DFY61YIlHJYQcR
lA2J1Jyp+HIypWd3LVg/gN7JiWz3vZzB7lmxsv+rhlBCLoX0AO5NE/IT0XRknSyN
L/bRp5ACZ5PB8pvAbZx0TM72HuFjzxbZEdvmIfIz7gNoURI8Dr2AgOYkjQAmVUMx
KuX50JGT5Jk+Y8ARaeAitzufAF92PasrF2b3m4BsF54MKO33orWu1cE9DVQ0GWoi
DXsrLxqSjp/rmTea9JXEeZm/7ua3pQhOE/bQwLFmyTJL282R1sFbu6A3LpsjQcyT
KbQXYCfZ8LZJKEIBY2nHB6h6lobOxitQlxoRSxQbDloowy09TAlv8hFbmkqlsPTG
/N7LRwQ3a7RM5jqP3OPpwJ7WBpZLDeKjWBIt2XAcCW6FyGZj4Is4Pc9CuFiejboN
yJLR67EY4EVp1+ho+surZ6FkGqJ0tCjJ5qiZcRSVXH8Tqcx1IAXvvSr4GinEb9Hw
Iv4UpjiDP8Ss9M/Ob373MdSI05ujBnra7QfCHNzry+yp6dTSszXfyVQB2nQitez9
jZyPd7SiAb90Wr+wiRr5obmVFTkVrBlHJK2aKmGBwThF7Hf3iXGKHZM1p13P5UbK
RSezpN6DV/h79DrWG7Mb4xDLUwyYKqDOp0CCKaA/A3CPHuczGPPp6wlwlq7tfMrN
pGhLeZhRf8hdWzSkWW1TkWVOnk6BlAANqh/Gs7twukyjX2MY9CcjYnZ0NT9vHKFw
VuruEoRHluw7UejKY65jzQg9L91dAktgQiiFHxApN7ywSZQ4xR0tHfp3SmdMjQCs
arT86/89ETtTzPOvC84Syqkq7MqC/EAr+xHe3k0nOPtSzLt3C21rPdpov8e5UhpZ
TIgTpyDRHkAmWueDOgqCRPKr9u4bt4gPRlY/muiYUXafJI0n2pAUz36GKTOHTpl0
ZOFDl/PK5lA9pNp2y83ouF3j4QL0pNagDjJrFEhfJl9qzUIcZ8jvzl7wIasTmpRo
2gRjM2mnhyUdoBxEgdiQ3ZpTjtt8yT8GJ0u4SoC8+t4IIS6dhtrzdtS233EmJKUF
KRVEtHVObQRkbbs/8OxJzQdhrGADd0gWTUwxtdLtrfA1JyMJOCNWyowAmLvuDezh
vQsl0QyYti4GEf0QwoolcyZVo93LtSPyOr6aqX+Asa02CgT99GzdzcuPDFUo7m0s
+RUJ2O7S8mqBsJcTJpSgATcmHA7MViR76vlRza2Iv3cwYYAmgUqNIjTmx0XOnjcy
braE5aUK3gyihNZTvaY+v1rVDE4b8ULVZeKeEKWMTLez+6C5MViKvg2cQhSD9x9n
9njmUTAiu60jZM4oFVV818JMuqzi4IL4FWMN6i8XgACfirBzpG+jD88HSpaiqPgI
H/JB2m2Yz6DJEB2vrnPkb+RzmGVuYpNoT9ArK62JfzFzepvVf05M6qV0LA4N6PRB
Y7D6Wxi43o1kwMaQfa8cTcTdZgf4q6FLE4xd+iD6+IB+WO8p+gy+WRTybn7RfRRm
WAl4d1qQsmLpxf1M1PXfPvvv0yv5cW5qu5pFxUGJ9ApU6kRfmpaowLD/nqVcfD1C
kSKCKIun3i/UVOrkeE9Zzljuwzzchty+eFRFhv0yYACjpDKRsQ2p/FLDDzWi3Af0
jHRxM97gsBPexZWtUDC9ko+HvYn02aCQS++EJtS1aIyHXSTwtcpnz6GC6snyIodx
cqqY5ifu48FrsJWw8DGANhCJciLxp463amOc8c4a8nw0C5FrbukuZJ6Vd+cubDPx
uMWiPnVHV8TpmgozVXOYOsvXfwruuIc+vivcYy2alfUUIRNYnCwiA0gsoo1AVAcq
h4CTIAyBqCdfWXFoc35kWmB+xMGRh4D48CxwXkOdXA11HlsoXQtWAGkqv/5hQodr
/VDs+2bXQWDF2n/usMgK9gka1QiXpUI601Q+KI9ILQ9RhQO3mvTqQZBi1mem7cXs
gSuHJ/j1hx49/WEDXzXWYxqbC0erekGD7lyNns5pPZ+i7a2NFEZ0PO+OrQCHTh9l
t9X7ZsgeEGoQ1kxCwkED+zUuLmwXIz/8Lixyx+/gIVv0BYtMs24Gl9Mkz9DWbMYR
BGAPCH3F5c+v2r3QXUxtaNbZAKySd7F/YM9akV9FnjX/2liqWdmJstmlADiHvaPN
traZu86ZNVf5VwFRgxMxRTWfPB7WUW4qaFrD5L4I3P4I4jIn23rtAOxQ2Abbb9V7
j3nGibrHWqaBbGu8HKlou/TLjKoNaONvipIh3v+ogtxAZhB2x/pT5FdbpQiYsLNN
cpUG3e0A3gfBL/r23N/ks95ByDlQEOZWelofFZvNuXIQqGwJjT40hUlCiH64TQg4
8RXBtqupsUJDLIDGrg0goRYXOXcY4NsYBq4JCw+Ap77pZbwhPMtaIVR/IU+zkqD8
KvX82Kp6/oZTCE2LZIZLhFVXXG8Fn03q25AMh9Dd/k9IN+OO02lyb+YufwHpT+pN
o9EpNaUFtCU1nrNocu/9ea7drC1SycFLGQ8vuO6X4ixs8h0d9g6FLSicJf5g/vg3
D4BOvf1a4FNnEmpkzWJ3c/YYvCI3dIsgcpq/UahTMYyO18B9usGUzi6twsQ8pPpO
LZqmdB7IiYcaMRqmk1qz6QBBiQtG8mIQ6fHcpV33Op9t9PjUB4z6SpqsL6OJkBw1
bwOaaW9s1qlZLCjmEG7J6RuLwOY9nz+KJHaJmg5Lx0kBYWQxOX5A/DECtpu/rdbn
FdhEQ2LiNOoiC4IhyonZ2xdZF9L1yvcfz633eLDeUg9r3gifxXQc3Zdugub3PsAZ
gql1aR/Vxt0pf7BeIgsCTfMlMa6nDzPtdFbk66c0XhAJ82Dw9l59yO29urjo82RN
UsLZ7gvrY97khJQWYzN0b61IJM+7l/aE5Kqk5dh8HCPUQm8Rv7+8dZd+J+aRQG3E
ZdDmvDe35oCsXtnOn6Y0Xl+uBOcIWcaiqqYEW3j9pGYNYOVuBISA0FAUxA6Whilf
zhTu7eHDV3/YAkl95tDuteMs39ROZN7rtcTb6ZcB4HtiISZG/0TwZfXaZX+p0/d0
YoW2GBf/QYi9YKuoV9VBCDGI0H76UNPijGZswHsiLU1wYhTkR5bokkzC4HFMzFcV
OPCiR6Th8CfRdabNdPglwKbR1qp0i10y6uD0anzKkn8h8Ij9vtFKsJcqfVhA/Rim
aewZHQzIM7+5YVRyP6bu8iQgFSfYKlf5g6ZDstXTDjVKEsOiFIKUxwaPsIe8ZT5v
tC/mjNd6Ocrni4CDmKMl4mZwnGGU8BCzU0YRz2hKDHQCIaOd/muqaEm/uBdkHDFI
cvi2LKlk/nw0Ahi8wUUpV6uVL43Q0ojdzOymV8KVnJ801UztRxA5XbA7haQsxfzA
wNkgjQPPmPJC98x32ao7vk1bALlQ+Ji1P4Rs+uZ8sr2to5Sw4EXlIAea9pST+HXl
vQy8G51v+jzGW0fI+TQVOgvqC7HL08rHWSnTFlcz2u7hStJm7Wg9+5bjmXs4RP0y
Od1n14j1OTf0+ar9LiqGMh/3Nq7cW4O1z4lajLbMTXxwx/2xHEa6NYbEBmBdR4cc
n6K6Dca+KKoOOlxF+2cBiAQwaChLBZjrvTsVJO//zUHDWUlTBAM7MocqVJIRAT0V
8Cki9oPER7rN7DY1eHGarU8JuJ76fPorn/uOQcUo0Ur8CmJn16q2l2RCvR2UGt0k
GyAn1paI8UsUHNTwZt6Zl0+T9iWOzKMy+dJ1NYwxvIA7ySW4gkg1k9+SHg8qO8GN
ULOPp6UOKEqf+NR53aRCmCo82+LDCA9V1gBIxLjuDoQ6IM2e+XjSsLMFAAV/sGR/
S75lwifdPYXd/LfBzbcvyyuNfMtOPeRlFOcUb2ZMX7CVZHEDRzdA5nrLcmBiruRa
11VmYbydgZ9APzPquXzkKR4dmwLCyTNzgNpLu8vw4/GwWhZODA6RB7TJQ5wQ9mPa
FJzm4VRgqHt/hoGgRWOBs1ETrUaawhhHDlpL/B5CX47f38+yOlxFhMUykWs7QK8m
l4h7NooQA6CnNChEfhayfGT1Xtkv9xSVgxfJXS8qab3ed57pSkeF4vTeo781CKjp
M7D6BN4+K8Tjynq0PC+xenpENuBUQ3tSFBqHLIWHXLzmUc1t2LpVgMegmtlKuNCH
dcZhN6+LgrxCgXveCEhbGne5MrMqzqVq/l46alx7hVKTZlPuuhIks4lvW5AW+aeW
bvzjffgg9oLX9HUacdfz5YQNs6ciHnMCi0caJvX+QoE0qxvmg6z4CDJpfXsAhu6G
Rr/HP9K51DuEw/LdQpD3sqeC2sFqCO/o9djpQSlDmYnyZr+0HzYT1gAeQgEpyv2q
2u9ju0bbD6FywtzLJZVUinKn8re+NKufyvAzsdnnLSyL20Id1qLiQe1Nb8x48rTk
pbLNqxptFDz8V11otuFzPdm2U75cOSXcLZo/uM9XF0CZsQOWL5PAM3Qj4ewC+Mke
IZol4IZxhtq4VOalSSSfA7VJDsZYm8iCkNvHQL3TsdO7zPxtypxQ5yiEfEwRLsvx
cR6YBLCguRDuitEi4YfgyuKDH6C8wNPZWQRViPBD0R+g+dqET7MjHL5wFM6TlCw4
zhVUgfCYEvD4v5jBteNxhDhUXupPgdt9osbV15Pxy3C47L3pxIdFzaUyC0sC+0yw
BHnQpzmnICAqHwRjJCUUu/rIh7a+anZOyiBsgMIaXNPjdbM/svICl/j9VXpuqRwW
ACzKl7Nm/ic3wUfBt6EhHpU4d4CMmV3W0O6xagp9NF+MJbE3rdEzhCFiYCG+8ejL
WWOJfGOxi4MI0UXY0O+tEwDjr4AZEriCUNEb6eZPMBt3/UCHeMTr19SdKz37Ptwb
gXuRXz7krZ51QM9E6lgoAuhT/puTYX7h2OivBBw4jmnIIEsRsBYqDzu71eNx57Ht
H3iKayM/xJhRNT+bmneewcR+V+9jIbtY74QcMVME04U30aMoc7XkpYtLGpowjESi
AGV0vWghpS2CFOYsiFHtQ+JoPUdKrLC4wNBDZz/MnZtJe94uSCYMTATnGu6K8o/K
I62DK4xr0cJCf+lzAj9VKi1eB9Qs4MMWS+wJdIUMY12qPJUXH2DRaU2Cg9wwdE/J
z4rr3cNDFU7CoWxTABcleJet+e/23Pgq/ckDuOH8/Y/OUAOaGmI344dtvNJyfvVE
HIQEkuVqBOwUJ1O0PyZwem6CdOgpNf06eG/JDHiuP6vkv5x/PPnR0zrS6l6O/CYt
qTX/fGEHmAQjsoKuifyC2l+YrrkAF5NSZyPeOOlTtfcgtQ1fkrHJwN1kSChcyh9N
8o8k+h+AzPiYqzpvMpa7KyOyNVU35u8gWoMbtrzO3F2olKWn5hFB7IMILZczCGAX
pmMmWyMf57LybUQdqFhV5VfSKAkC7PfEgvTyIr0LahV7uir3BhNxbLyEoLLP0tyq
lfg3HVAARRKQFuOECIPWZp0Ip42SAfgc0/jjCP1OTsJAub84NA8iffaW4XQZ2t+7
/FOAbzrSQT8RLeP/B2SeXSRTV6e9vPhehg8Ak3L7ktpcT2RdXe7TojQiN7v9o8pZ
yprfkuEIJ1ybHNR+8/vUDYFUEFRphK8gpt5fYAt9TWPUm+fxr8EHiw7VVoejWxIe
JSrgfpPtcIYxkZVcVDEJ6UPQfRxvRDR9HGUeekr7VygNF1TzWKOTDNrW8zg6E05T
gdJVYh/hYu4run+kGiB973GuZ6zcBVRy5dGi2+u4rwLi3ImM3ERUNtHLNwQKUEs2
euK8Ny5Ia+fzHX+s0hL362Jupip2ZfwN5tCG2qafWA7I8ZSONbK52hf0916pWQbP
0YGNGv34rdHIU5xhpIlWGaKVNSQ0/pibVgkibGTqWS19yoG0X9vjv/SeTASDBKB8
IAEp5V5hIaGHUXxGVkb7v2QIZFZUssQ9KCxSRGGIUac1TTIBeOKTfiIaDHW8a/fA
DMVB3bMBO3aINma/w2TU21iJDr31QSlzdjTE06yBPgkj7/1zJ13E+zoiWIfSTFiw
zB9PzNn18CoTHGqpWMVLS+iPIbmKYP7o0Ag9hY3+9GP2BUMA+LqYDi1LUU38Op++
9qIuLI+lbXEaPDeCQJXtTRwJwsv7OTxhEcarRanoN6Sd/ZDYSCAThgk/dZ4M3Aph
u/KO+2qvFZnOFtRTaQcTerW7faHl3yIApePXzuidr8khv1eY3XMQgDT3RQHIZUqL
4Lzbkx+HK2SgPHQdkTZwxPooE5gwS8f6SualsHy37FhYl4F02ZEYaGwaHc4OhqXn
lYHUUfP0DdmaDfgb6zC5HtCoK1wK0pcX7Exr4RlJyiVoNqkqcrYJ5njG6XHMb7Tb
j4VWEBxK7l3B8keWxiG7JOEpXZ9WYjd4v+cx94/ZW/B9Rf2+aN89DJJcmV8SbfSG
XW5hT8kr/e6rMFkFrjhAB4NUSoF21VR8yEOm+c1KGld24tzKPAJXmRa2fp5faB0f
/egjx6HZy1T/mcCKC6YQmTKZuFzMBd2uU6/k73xsJA69ogv1XdodZNtqfXRuxN6s
liraF8mUGh7bh7jTmL2FENCy8L2lcq6wr7UaerZKsSieeRTYnp2fRfG86L9eKXrU
HlZtsEXEec+QF3q3RuMSiOSUr+JQYP17TlMTF0CayactpVZFES54QXf7UwnSfpgx
y3OWhBBt1RBNL9r9zz6cR8No4BbZYupj3xw3SodxTqxYtpknaFo3NoxmfdK4lL8Z
4teC5IcUhmUeLj6XZ5frQLtGgRKH6JNSxZdEuEdPxGXcNTEN+Pjxsxm2f4n47r2Y
c6WY7FknOVvobo+YCPOOdJRRbc3fMWCu1f5umQmqsjVjxYjm5+zIqM2h2cMFpH5X
bSyw20bbJtFRDucdrvRodIwurA6peDkTB1HshcKZ75be5O//YbodK8yjZucrSzHX
7lAiCANoGCpvtutjwtsXVe9Yu+0hoJda+JEmdhtVhskb+O/MsR796c1VBQwOchWt
S8L73IzMgk5sLhf4UubXrJ3wiMTfXH0nTsY1Yw1XVBRf1h8U2udADdnfbOQldUZq
+PLBYaE7dsu0xnl5X4jNz/OCxGJCVGnG+eLSd/dxrXTBwEDUg0ruUaJQvfZhgbJi
vaOkZCoRtAN4hEXlrx8v90/LHUcKKc+qLWB3bPRWbzz0jQr4c5zH+BpqE+CQWF5n
N19315D5FDLcMwsjy8L8OP/VH23HJa3nt9jzhm4TT0DUgATXZBY0I8Yvd+9pKGTP
Rl1cSdnWgMzbbhKnmpDJJG2RxEAOaq0Rk9UILwxgFi5T8lgiiE+wSApFFzM5h80w
v93Oz3DpPv4DpO7zzSUzmDvL5I2EtK2IcIJbVtdkVGdUSNlT6Ovbyeclf139RmCf
TyJ16b/ZNc0B8POHC2swnrzHvrdblfG0rT5KLy82OpvVyqe5ekODVQmiNcjzGnJX
7a+qmzdCHtIQoRpqpEroHM5XeW8jE08Bo46mDwGK8AAlkmFsJmbNwVQtI6prtmDF
2XfthOpfa5A3ceC2q61o0Vo97OGJkseEozDxoforP1dSN/MtOWA60DLDRAJdSkcv
VhzpIYU4UqWz2LijgpfMNn8b2j0KJadUKDHMwws0rt4+epzxqlRq+JF/idsl7TLK
uc9ntSMu9skyy3EWxQu3+Y4UV0G9vKE5f4VGkMQOWTDOpiEe5Z2D7F9Q+xdRnNJ8
69JKC/loGDdmtf+tgxOHG9SJ7vYN2epxRn3IX4XWQMMaRo33hTTdCGfZPBuF6zj2
M4TS4hvKWqpt1QJNfTg63vLkoQi4S2p+/c9HkYtq/sr3g+jSlqKtU3Qaj14+jz3j
EbH69ZYJSIeHFP1jPRuFZBYqCsKbTMMQ8IUdO9sbfrNOU+jd6+fw311nrtYjjxY9
j5uKeznkg0oZ2eEr6cpQUJeogof4HbiD+hqT8Y4cEQFEGjIquO+NO6dIohs6pgJj
4gyQbc0Dwh1w4rHE2fA/SD1CxsivIK+Ai9IbIxwi4Lxv34dV97rma90pQ3GGM0hz
4YYqv9o9Q3BNM18Gg0ZyY1fOwXKtAoj7C8O53Jr+TDisJsKxFzvEVcgWecLSj/DY
aFzPW8zttmnW+224OqwcobVK/dmYjJSa+QaslMu1M3CyIE/7UAm8kHnL+gPj8jit
ohH+kYy00PtMc9iTF1uAEHb5x/aN7R8N7bPHelKi1ifuyLaBb/xYm9zJ/+7jh9Ls
dILOQBpSL5h16mVyRj10bibjjyboIa84Hj/YQVXuPQFYu6ABJROv+L+ha8o7Tirt
mC4DLWhpwnFDzmWpF1f3u+ynC25jGH0N1ln7TQUbbT4bsxq7WyBfN4owGnC/A5SJ
VdyNQoyzFP9ygbzqHLpDMVv3j/SVbF6AqS4WUUSj5+y+qRZN+sg6wSCmJtgsVP5K
ZDCPReAtPBRjPLFxZRm76HCoodCaVSvBZ7SssGhxrlrdNIemB+l6yuPHqeqEMg9R
ydNHZ85bG4BZ2RfH8wwjESA9XzzI9xTFzpXdDcl7McLghDCM7cYoG5CP5yxDRreV
KY9fZFs/Uf/UMa16yVSL33hPU8+QLTShAyg+Srv0NARgrThOvb3pjhx/PN2Ls5o+
6nHSNRVUNBKiTQSpeIkeefSlIdCchtYZuSs3iQlxS9mW/klUoUEnIAhn59WVjzAV
x1wlJifDoJQtruWhsUA6c3K3yxwBRsoWXet/J1Z6iQzLbgOHOS2zm+6o3m9Cq+oV
OVA+ilWkYR5IOOUhURN//JUXz1byyVBFmkJfRmEOWUWEbWb/9e1rhwhAgLI2RqYc
HhweYY7RjOzc3k5cDjVUsHGn7et6CXsC2sqRR3mCvwsRzU83EhkcQJO+9XwjVooJ
j6IxZZVdzI9dS5+O/Jf74AA0lFVJRlZ9HvgqK2553k10iLJ2VEctfsfoj5v9syah
6v/SLmXqpbDY+Ykqd6/EE4zyjdbhsiwJiXBL+Gm/A26np6Aj3vl85E5tJzr8B8Oq
24VlvYQuT/3qMJUKzUnBbIPEFCQurQ0aKwQRYuUeMH045cBzh7ufr3HDCpDGWrDm
R5WGut2cJEeLCsKeYLaojfyN0NqD8fjGuT3gcFPtIPUOjn0z7Lr1xs9ZJnIcQsya
iVspRkmvqeREWSSCmi3Ka4Zqglw0gOj8MoksB/ZKbduqshE1TfcVFvXi907u6ZEH
RhjM6UcVfZilu7nhMpB4WriLaJm98dTdP4K5l+uE6/GRR7Tx+/84hl7V1j4AkjX7
9ShZ02k1bep7EbB+QS56GBulgfMQ2aHJON4Qo3roTk4zQ/arMrJdm7Moa9DfiSPR
o1bihfbE9aLQuAY06uDwmArZ95npSwRzHLXfu+6olkK2IrGjXiwqUGcjnNICMnc5
N67lVTi8Od95iP5UOKz9eomkQgN5Us86r7j1uKoUSblr1IupRPtEGhJvfaXafl9b
Mo5obXxhb4z6DpCqwWCXDDJVbu3H4PdGu13CSLC38GoYEenie+GxAQpuRKkpIOdi
oEC65YAvtxpK2HrOevro8vkoJHoL1xcXdRpiPsju/SBAg2dQ2VjvrpDafp7zQ8q4
bvWRcP8UWPG2r8APSQiJiqfaScl7xbw9jMSjKXyGBJhdTyuXCqnQf4Ymgc8Wj8Ln
sdzlSxAQsNUJ2epzChqe47RHi1EZMMhTDhTw4z9Udg5iZ7ZecTK5dZe+dxFdw0Jv
ygvLFbVb1Ee9chH4jUurj99/BaCCs2zHUaPCEcofSxaelpzv/6fYP78saGuAmI0P
2fRq0lfsvwt5iNyAeIUIh/IKT1ujzlPX7hjEpszZSf8iGL7QImnp1tjZ3iwqMHoj
d7iipMQopzXQeo2BzdjUGADIkH60C0fzAoksXMycgegSfieP9BHTsSUBJmfhvc81
naDNhu/RZIDIctzHW8QkrkPP4wtN6WpY/yx0T4ZrUdG1ScPCVTrlYTC/tvkeafdP
9lFJniVn9yi5Uoumuskc8VeH2VJQbpPt/dpUK6KBmpcsVla1x9rW8Ksmak5j8c3g
yio9nJSntWKaNvLklfrO724j64U4o/Rarexb97e+/4Jt0hmOCOPvUkvwE62aICsB
tmRZ0+j5PjZwZ0q2IFezb2FyrEBwN3gYNv5zdi7JS6ayu3ADPHh9VJBcOBZOjOeX
f0b8b1slvfZJ8F7yMn2HNPfMh7DfQ6PdecDnX4ZELOloSTUxqbUwS8KZiyUkBpuW
eRUmFVEEIEqpzo7bUVRk/oBXQpbW17SA9xtC6NxILh/t4/vqICA7xrMsl2I8jL4J
iJ/1bInssYTto+KIuM3KL1J/lMm6VovPIz4wlhBEwBVLpAZy45hHwgQJbjJkd58e
CNEFyYinclHvJhXUbgxY1E3V+tOt91Ew2keaZjZCFtYDDSasB08k2KFDwZj/r5x0
IwI0RdmVoKZ0VeE1p/g/n14DhtAXtD/cnvs7xihIacFzwoPOg2xsv6GXYAfq9Bm+
bxrKi0IbnO3e+sP1Ec+RMWMdBTGVzXuMPXMn5viabsJ4ss6o7iHNKxhxlRECbDw4
Ce1xM/oXo7VZ6iIvH6f10M4ue0WoD9VlTzXP6FlPERBcUUs+x4LBJAJ0qGfZl3ij
mN3fZ3Yhu3ZA0Xw2RQz/19CJFPJttzbqFGZZHVOnrES09pOHzqxMMtAr+ElVxbDQ
fqlMuWNCw5G9KLegiFCk/k8GN5Z/Q5ttzEkke+3DPyipisqvsnIT2dUpcgx78rbv
xTLcSAisRDyixh5OAuUNi4woLZegHtZ1y940geBcYHUul2HCdsSaCgXxCXf4z0Fs
2jRz1+qWRw8GpSK1/S5Q4myNxQEW3XTDePfMoT5TZYvZg/x0ALt8NOAx2cfK+asR
oCKlykCmWIXc1uiItQPWfo9EWQSQnwOLapWYg2rJs7goFOveK19X7FrbuOR0G0J7
TvZL14RebDBI4GxNT0slwmpV5m37Cwmsyarf2a9Rc4tkhbWq2d6EkXohawEhwCQz
YluLVLBfH10utrdAhE4g7+Sx7yRQ1GOjhfXHBw9iF8xZ9IL8M4Q8Qq4jPAC7dSiL
F8D23gCBZqXe2r0nCicqAKXiNXi823Yn/WICX8VKqPrd/x+Dzt/fAfOL1KNYeTVH
D15lm1j4A5z//dHgN3NCszRmNPZI0dCLqYyw8DbCScI84VvZFidULvAyqbdcgk10
68/6l5E/PRjuCsbz94vB+Rrws2yShIN2YHhh0aI7Nttd8nYX1x0fRyTP4Aq6886L
94aKL0+xaZY8hlA2POMceoe7OcQ2EMfJEAcZVbphSzJk2fwT4LIfHPuvpc2FZzS2
ZZxlvtASW7hxzgIS3eyOKNjP3JOJAUpKniFe/WXwxYoZA9j03luTMSTSElOJZUqB
ExlynWmch1Gz9o5Bp0C2PQqJ71jBuVW8HPY3qotooR88XNDWViqHAEhbJ+c8nDAT
QPda9FqK/4lHkEHG92B7ZKjS0veppz6/mChiqELhSW43dNfUd9nXTcsE6K+AkpUF
8TJsNNV/+U0tgiKwRBwGgNbQmLePtWuPgKxfTRtW/Li1juyGfdJGYjkDolzoQ0kJ
P88Jzl19gAjK0S7RP5+Z7lubtEsKSw4zKvYWOJns6VzDvYQWTXEv3jt79hJOLerr
k2c1MoQInt2Syyv8dau0TMtTaYGDX3zGmBHv5a4NdVIKX0Wv4Z0ZOja96iWOf2m0
d3r8FLm1Zevckgn/mLP/YzKrNoW8aaJheNLRui1/tr8eal5N3V+VH3eos7Zm08By
GFVna73KUbEb6jm1LZ8djo/Wahwgd4KL1QduWOeB4DqcrIriQ8RAfPi/OkcDOzjM
yrr+Co0p2F8LnvBt02wdt3+av50CDKXuVdMnQW7exXo2KQpc23eWqlUkHGe3omVg
wwQ7oFoBLbGImwW1w0sJ/vZ9fb1Mg1XrYNFmZT+P3ClFAT0LGuZCGUrGJSQMQa+4
jklx3bhJvjWrGk6OAohry3Sxi+RgiKRt5t0qsPQRkaf4QtsKi2yqzokklCF4Rctu
dABYhFIYlzUu3dAI5B+243VL/88umKr+nxzxUi/f2JHdHaUcH1mrHC6G0lVXxxjm
9vUhzrgjmAHhixfyINipBWk30oMn/KEIpm8CAQSyfJetNk8veL5nG9s9f7JINOjB
Ov+8KQJXfeFbtBPDkuYQ9b6W1kgMP6sMdvZ89GL4h5LATP8mnRpYSBngor9nTSm8
zg37gScq/I3cMAqVPJj82QOUnYOHfzkLcSg1HefPWlEEU7ILPpG/T9yjrfTJorsb
gthqKhny47YwL/8TCY3+oRGSvpXnXdzWLKTKPdZnoOsSCLQr/RZT5wS+CM/olExr
+sUCaQCmF2PGu36nLpHYVremQDnPhUsL6MoVozcmL0IYbouxdvDRvxBR1LZOIEyn
f+qzEVE5H6IRwXe0RjCPKfSUWHou5BWu6PPPoUKqfgVD+AOVVjvvMPRgp9BCVsph
TboRaAI3kIgqZA4mWAiBYyUINHMXnhUFeax4avC9vX2vawzaB+DnSCF+Inhp2Fk0
YYXmql0Ht+fEN52AJ26vUWx8HJky/eAPadGzTvOaxD3Y1rhXBHpumZs6bf95M2U2
EVR0o8h+vV5DVlHuY2Si6mVJP97iclvox+d8d4VW+Bc93+szCHnapYz/Y77/cln/
PbuOIDccjMU1RXpfQ0KuuzjU72/PCHMg2jg4a55UVhFKtcMUwb01h5Sh0iMVEtrv
hZ6HNjzJr5Tew0PNhilyaYiVTHjHfrZHm2x7Wd/RqHFjR3FPvqEpgoXx2aVjsVSE
BmfeyjI+1noh76TKYQpDQIUoGuska0j/ebFaj/HJlOJVZG+iGTBH3eig27BcEh0m
Stx8w7KLnLyv0OBF5kyAwp+EDyjKmzrvYX+0i/XfEMA208K4Njtr3hq00ALEvUrM
jML9WfwpIUQQNT2NVp8Tu/CA6O7I2nKCMcNJ1RVZ1rNyM4xOZn1YnzhLCVO2qj+z
FPxakzLEdiq1v7NLbgiBo9B/jMvegWtiiNZ2ZKOn9eA7GtIbNp+rNNMNbHnqZWvM
yT15UtbIR6NmVE32X3TWsW650/XY5F+La5gLm1jO9eNAQxRKD63Gr++NXluawCqX
f8IA/1/hnjtISTd4wMPcGwkys4rzTBFUxRdBrKqFEpn4DBPzuic4X9GqkSy8pPb+
fcoQcmW8gHyjmo4bEpIs6qn5ZCCIHbQIEwRQ1EbYA7SoIUrufntqdMGPG7kgyl/F
lfkpCWtNOXnH5gCY0k9qaMuV397yUJJapnBdCjObWcrq1RCfk9H3RlGS6CXvzoRf
Q7Rz+uMZsjEEOSC0y5futkGigmrOiPRFbpEutdSI42Wb+GYfDYFfao9l7UZDXdmi
sk2yyiLxHbXZfUz2WqhGH+g4yDVqNgThKSbMnYhtpowU/eR2QpZOrs2K38eZxD+8
6vIozPfuVOI1rJaQG0zGIlOf54NYDYJdifVuRJe+Tog6oV+vl2EKqPy+QzdhlqOY
SkTPmxXaeTRcMjD567SFFfm+NBqzGNZ5irbOqV37pJlSfL47I78N5bKqCxEfWu5u
1Z16CUw8cTbAjU/YHVElyHgiAGUXNkQb5an6By7XlcD6L8QB+UlDFnorRwKlYBkC
zymyBiHaZ9C7OJmwmyF3hMKGDBAvlij24tNVCYl3SGTuZhIHRLXJmUwYGkXoRXVd
3KpR5LxJkqpv4do4sZ7+k9VLU7tJRzzqea3TOjxA3grRYuBc6q2yga6fnDQTbm3O
uDQyCDJGqYmOzxVc881SwzKUHhZKmXZbobro9SEKsgTTVSadQq+0cYM6HjygG9Au
rxxzoBmz48hfBeXhLoOHSx6FewkEa1Zl7csKBkTMLrmuYf3uIapmFHZLfW6N725A
C7e2ycGtc033RJxyUXR33vhhMTLWHM9H8kHeXGWXVXRmX07ZzTER8HaUOswNk4by
xmzPmJTCDUh+q8Zmslr+tJ3JC4llz8w6Jgde25JmKcE+o1eTnirTX7NHgjp7M+do
8eqIdGhj8pElPdkfdOGmxojpkH0wjKAgflpHn2vv38dxt3fuuQE8mEH1YHFwAvKw
ZWF6Lk4NhyODH2wEdyO2lyaxNdSp9mQr4OCI/i5yU2fBfZP8+U6l4ppHSgjVWhWg
7cq2j/BoJ3mRyQDs7C1ysBjHmLdOMUZ7oCR3keOcksgCf/4wVX0xx/NMGLZBHy1a
PKn3gDoQ/4jKI8xesjnN4JKRouW/eTq089uN8g4jn/m77MzVD56uJLiWefPv8ixZ
AgSgl/cGQzx40VJkdmbkeTGknccJRLfy5JPSOBAxxszzcdD6JBrpxHobQGBEibg9
qkZDrVne5ZCb0Zi/UVeXv972wV8CoMJRB3hhyNL48aE00OfaR2TlYMazgMfycr9Z
mrwdV/jcu2Q5jeZo7NwGgCazh+ROhmr2kzvk7LkFRalJiAL9Cs+JlmcV3da2CUak
T81r4H21fg+uP0X+0Mp4kCa4+ogYkpLaePj6exGfgLL2/YTEYAbcF5Yag1EZX0W9
xEcE4t3jEAE6z2a1Eh4PROFUipQ84oCkOYpMzH3Scr1FUmfB1N+iy0BhXHIzA0mM
ZiY+3ekCSbweKMsgNMnbMIagwkeOZOpi9GZ5Q92JYAMA8Gc4gAuo1caf8GUo3xx+
ln9hKUpQm9atjjSIiPo31jXTHKKJ+ODoTa7EUkWDPnuXR9j+lbUMeu9qLKjcv/6/
uSYwm65ClN1NFttegCw7ssq2VdkLvJTRTP+IacgQVm+FUvjN2ExP0NXL2YvlXE3g
X418LUPTANrn3/0GsaI7vArYaCPBT5MI5CAaJQwmUeev/Wh6pIOOLcqKaGXs0J6x
yom8xUerGEacylgCUOyPaus0ImynutLXqOgTK6lPNX9UC+/DbHJYPOUrsBRidcPp
VdBHM/VlbVU2dH2/dUBax/XhNSNvw+3p7E4ShO/+0nBJr9eBuXS9kBUV8PzLjmM4
JbkIY3FuEl1eWZ5c2xGR3/8Kb4qmnD9W63yBFT+TpbOXfBZwFHkppUyN0tGSuCrl
+jpVP1zzB9JHhIooPj4gsqlKDK31JMyoVNDiNC0PzYOt+mxQCERuJHTxRypH0F7Z
qTmknNlEphlq8v7tIDF+rmyaJvugjnRavfBJ5qJEyyyCO526BbWcQVuU17u9bq9R
xxViwLG7z/2OpkQlg5U/OotTcB52z3CpbsAh5SXTQdXUKVFivZqdJx4n7Hc0f05g
FZY8HdSyY/H1muWvZpx0o5lERi7TwWZPeo5vft5MZPJdPpsf527xJWJ0VyfHyzxl
dBz222+e9z63gZro2kl8UV2suUVHam7Y1bE257dh3sbeocFPMdL1zQ3CL3bhgPCq
UYbOvYky6wBJhuLs/+rl6DX5aIQcRKCkRrPf2afRs/ny9cGlbLa6QCG5GUN3/1yU
k25xQI6JW3pgNLPKwNLAqrNbGqNekO1chUv5iYZ0quUpWeEDtLe4ZjKCV9OsfZ2c
1SE9yjEB/qY5GObpi1y+clPTivezDv6r9Y7mvsMEP0EQW388UOlTBiAdTilCQAZr
koT+7NcdaG9Itu2H/h/RFQ/QRSlMVZsUPEgXzbJg0wlbtEKXbfVlIOQxA7dCVgJN
tfv7kRaLfcVrHyTa+/wMyVWXo4ph+iNoxs2PCmhw1NLL8sacByhkIVj6GOyRMfPu
beIFjx9OwDM9kiQ4qZthRuKCtGKalv8+GTfHqkET4oBMUGI6lgc7gHkvl2rS4ED2
FygAcyTk1Zql1UXSpi0AnjSm/ee5rdmYl3rTaeQ4mSaL2qtjQxFrPv9VY7FyuGII
1eNSy1FI7roKzeAx19loLA49r0wtwVKeoyo4NMIgzmNN4W9e2DtQ2dWvoIfQPkJU
Mg5UTPxJfAh07/eQkLrsMb3U3pqvLmUVjBkzWYte6RwJQQSUT34rAsIOmGgWc0lo
/H66Ji2ystNBBuIrxjouPd0mXa63AkH5r/LnTmA+YqNZBvSrvQM3GkQjbptQ4tBH
zxq4SU5rTiaEU7b+eqnmmDwHuxOQN39APUsEZpFl7EoSF09Z8Beg4/PlN34pN/iy
u5snSx1/NO0/mLXhT0tLvPI6UTRR0XuTg86HMljJYirqHRpEnFLDzNCdO2e5+24l
5BM+Sn0vguONGHYQ66x30UmdpAnw8whvUj0ahuIRuGp0r+c6WzdyYnYiWUofIhk4
4H4xx4wEmzeorK1MKDE6yiVLRiPLiyhqHsYYkiyBbH5QqkKvH9/BwFxxcw5RbpgK
NdnZA3981aKq/vG0iadTUM150Wj4KUelOZF3FM5whxa1cGeCOTYwIr6VCTAa2+GW
0j/CkFm57HPJVWpFgeCQGlRX5ARDCD8v1dNVdy+QhfGaZJQEFXxtnnPbyI66+nsi
AS1BgmeSBRtajak+0gzOWU07GVjQu6La+tAvx1MYrXM6L4vARecSbsESwWTSLBlR
yc3/H5GIUvfFNjz6vZEL8nk/E7dpG5Qs6MN4jzeftzIp8eleWVM89t+V5vczNaWT
EGc2pJBdO2sKbzHFlV+A5qhVZLuXs1jWwMZC4siVGMcHx2zOJlV3SfhFQbeb2Jgy
tAUDFwVhQG85YqZSN0NvfTXyJPymGLJo1XiRTeylRjtnp02h86Jm/GAMODRaGL4s
OgZsuqkvYnMoTGTXn++Ns+tTHUjl47u+ffGuOv3l3shP1JHKZ/OoSlXhlblZKxsS
qQ92P7XTklpnwVyV4st0Ku4i6FgWBnrHhT00BmwuRUPU/WdYeBRS8SByS53Zt2Sj
mg+vm2ReS9iqKMOxo7RjFzm57u5RSJvtUUINmZC6NUFbmo20H7bPkGr9ldmQDjQU
zGVH6Xfk3InqEOn+BAnAXE0+EOk9chpuuQN/jU1jqNJ9HLRrXimNA7ZBc0Yk8jD6
ekX6kxgmJ09JtOsD0OOn4GkCnXZbLlOLehkfENHBrVklHEDWZ1d5p1GZvGd+D2kj
8ol5ZFguOc0EZzOUZqDKSiWZTuuQ9j+ecIsJQhVaunuHpEdZEeb8ecQgGk5R1fes
iMb98Ev7sq0G52F0U//Tcb9ShY9erbiMPKCN0H01vs6bBSAUDrCihkWwdiryPWfk
T88+hOp+FolZlOwy5PAkOw/yI7YV6HTH50byKNpiM9x6r0UD4pzDhA+GqM1pIyfr
wvdN0k/Qy4jlfq6iZVpUGCAqQ6IdP04JMBZcH2axcFrbrdvZwkxhCCppDewhFgdW
8fz9euiOQ8PxnnIXuUXORX3iyUth313bOoiYfqdWV0ZRWU5yQaxFI/ftn3SwTo+E
aSYHr2vsLSJbgljzPf9Wfixpt5LebZOlt3QvnLv1eUNkloiC7WYMhYNIDQUOJ1yc
AJgB52UR2P2EjxqKSS5GjqYiG6kOR+NMQbL1JadkWuopBr2B6MPUGP1D8PfcHaQN
+smM775YGOpXghKperQwx/qDF+fgH3FKumsUFlbGsNs4fGlNecsTMCh4REWwIf6H
ThxwR04aHDCYA9Brx52WNt0SITnYlvSCuxmnbo0DTU3Tb5ZAfWs+1V0YXCGV75U5
NQSM8Z+TMGqgnevJNIb4odKy86JelCdPeg0xisuvPy+7qOw/tXw2fvD8c+1yA9Xz
abTpMDoGbH1Ie4IXlpPCjiLHAGIqz6PSixrXPyyZURpsnfe36alfVEDt31A/JbWk
QXqHzSWEGEsCZlDFkexwwgniCIK59SucuVk2g8BwKt7tSUv8+ONGkw7vg5O774ZH
PRTZsShSBYJ5P61H8XK4cj/m4U6HYsag57GfPq7EcdFKxRq0v0Xngu1vu5fDoiFQ
xHmhWw4JKK3oVdDd+IfYnlwxCHIDokRnw1ZkrR90Z83VC6OIDSiHmXGuUwLzRI+I
TqBqeUgdQ4dYKPaihqHa65+/1foDeS0/BbdssX1giOORK4MY2VbimAh2OAg4SP+4
Fy5rwEQzJJabSJPFKr2MfciKg1cEKIZK9Fbe/MLXBqF4cbVjdE1bw7kI2W834UwO
xJK/QIbz68ePzFQOw+cDX4WbFelxTF9gvxYABxEIRdOXFZYYh1APz8zf849Ofbxo
yRlIjEde2lRGSzcmGlfUccAlBh2RO5Fw6Ahm803bXpI3FrAXdGPpNgY1d8ZEczJK
alJ7u9et9Y6BuoKdQASKzC81wVrUXlY0iQ6mFDLyKdGHqtw+ljJzdPYMG4Q+pGhE
IvgefbyJrEFkCTfJM4OOpyiQo/b2ujEnfEzcH9vgadVdpYdxkj/bXEwkIrt9wASX
BZeBWzNjWtP1G1rAvB1PS46ctkQrGL1pKrAe9UkpGXdzjnEKacjegOYDFxoOi4pM
dN41WoqzCzE3x4F9NQrHFk0JLt2xoDNLYVy9FKJohB92tBJf+3YBdvRS0Axbuczf
+s+e0bqipbuZ9Cik7E/pW9s8pJCUfPRZRz8ZKKMXu2ZcPnrR+L5rbZTE062zdbux
pmKgkb2t2z7abSwGZOK9xEf5XgzuHEDpr8uvqYM6gp8dZayePPr5ClgG1sXlvwtE
MOs2gXKZVtc8gkhOXcZ/O+zX+c21pP2Bdg9e0B3EzKtTrLeZH4nhFDBssjcHX9hh
IaYoo9GYnh8UKkuYXCJa8Mlgam3gxFYRy2YYHqHI8JfOwMgu50W3H22FN3WFuV5O
XkERQOz6Dhf+cxLxHawaYyVVtjCnrZ9ubtFAncL9jVKovQEnjjuFPLXDGjKyP+21
f78k/wlfvzKrBhvSvJtIDqvjtWk86yosHenNZqc+GoZcNHAaNS3lARhOH8yzKQsx
WSc369Q27Hv7FfLr6DnZ7BroJBvHHM8Pi5KTuCXgCbhjo2FYWFC37vstfHOCBlCB
7Qfk3nZttsij7RPARYPg62d/I5nOKtWTJ+7reD0cP60j90EIEHx/U0OpGCVdpW6M
DX5xceVg6540qk7FxUPU1fi58T8VyZLVPsiSaWvCTMGG+3D9G47awXs5/PiJSc0n
aYlAykkt+ru/N6rBCpVzvQMOqf8RcEAvCXw1ZgSz0wHWvb5T4mp9U487zPXH7Crc
krHg1AyYBVObMthJOrHPk411yZw6Lwc5WTHCNMLPJif4jpKv+MvUVpLstsykA6OJ
Y7l3zcj3nkL1aJUROBMkVKsDixVhh8rKLfqGqU+/N2dsYuD4AkzTv8gZcgyjk7fP
D0Kh0IoXNp7CxV6Voec37hEtSeNZ6/hao21eNtrq6wtoBLjcDM8LVVcd2wQnfAkl
sC4iVr8sje2oaCe5o/iahaHtJyAKTKH5z367KpB8AEIuJSWt2DGbjH3GeQZ7Esan
LRC7sLYHUsdp7hBgdyLSNnzkqr8xZoVpte+K9W2faQl0uhqPs62Ew0//TlxvtpIi
cMVTNc52wCIIPx5mxaxTUmw7N5xN1MVgxnljMKZkWTB8OfddY6e1TY2gT1S0DEWd
pZDMjfVwLG/9YigVVoT7niJYQ5uC3HwCyw9odWtmLrrcNx5U1rNsHjd9IPmHzX1W
STRnmsutzIlK36RO3mQY3Oym3QH76AgcHHjs2mjm5PTeHvCLgjef7518hqLrHb06
/QCoRSDln0LuCiZ3lyvLTydIaObcq1Xl9Y6V+9NbM+PJEmn5+J/FMSIr9vwtlvsw
9jZX1rOMm6YX3VETb1uBi7SYKg6wbFT394YD+wkFHDYiWsZfN05mPEwAEs1i9u34
rk2sE7TNFbW/ugFwaGlnUPDySHyXRsCcVU1IQFc2lhWnLKUiM4vJ006nZmZS2m93
p9fdh4J7V6RHIk1i5j5qnnGlYxbA7ayTC8b6D++ljAKlLtcPNqYBsngPmMRcS0lb
JwuwzX+dg1sPz8G3tue+xj/OvRAUjPKmn1F5IJYeRhO2vgQzLroz7TzwpZQAPHx+
sOsDWue3D7DJZtkcrNz8U9p+UD4kbd2gra40IYMKg+Y9dPW9lhTac9GFu3P0uDpB
04+UmkLyw5id6N4yg0GCynMoRY0Ue7DPzMDWJxuvmIPsPvSFMz/XJw93zjJ7bo/a
nBl1pTGOQzxVL1J1qm7x4473am1f5Jaxu6EjdnNxm7EmGot8HxMvSmsf5ozqJO2Q
I1OvnOaykoPnimZSDB5wqY1dztJtAgpyASBP3HhaPlwbX6Jb5yNexs4eyV2cjKlS
6KnC/OIzYjohPyVX0VPY4aSXNaB3uzksa/hxn/HowsHEpgNK0YnlrjeQZP4/zFyd
73CLMFQ5eniPSHkue/uCye5573ijnIa0F8v7wxGcprFmwm2/2V2GxSuYQd517gSL
9bUz9ol7DJiQff0QZlT3SFxWzXFshDfyxvRT8qGXezrWM27a/KRRUWsYiHnQSsrR
P8BDfy8JErkY758DxDZ+lsuqQmy09n+RIBAl+9MuiuC5puJZLWWNyv60izhN82zG
Rsl5w17dV6xxLf2oKjOBaG5umqJSvbQ26SQJSG+v+eJtNu/izmIwyTTGm5V7bHQ3
ZndDylYijyGnjA/0YXygUJg48kcQ7/S/2zUvkpU2s1ALqHH9qnpS3CG8/gxrEhU/
s5Gl1C2yuoOkCNwgyaAGcVYs/o5mQlug5neNaogr5Rjw54ZhFBYVMQrUOK4znIqo
0AbS8FduVbdbV1ErLeecAzEp66Wt7K7QxfkI4pSzuRk6drJxYvGgLMK+zGAMLv0O
3u2ue4jkSSF2ioGPk6tfJ0+qy/sFAh+34XYFM5zfAsCndgk0CwDn+W3UOozhBeyC
aBgTFONc/ClUCh2tJQlziSV5rr78TTo0Kry19a2kI9IcuXeT8lI5Xn+krq+V045J
J5Vk2zbFheD2E6CmDw0q3idB/cKo24f9pYPxbuj2mYWigDM2O41lwv5pxEnVJRnc
B/BrsD78czZ5FqYGaRB1SjEOGivR2vf+B1TKlBoA1GnwWmA7I1teA7YnRZfzEfk5
ZACjwf6jDL5PBU2OUOWsIiev4MQFqHPl9gWz6Uh0aXeMzU/P7+RSgp3ay8LXkLfR
7/EM1lqinaXUw2r7oaghNKX29sWrlnz/8kjYnvCYYR9Xhhl/WEkCrltfNB8eKf68
ezrph76tSKt2bhYyTByP7OGg0GPstAjc6Zwkeq9El0lf72XQy4XYJpd4aRNtWKVh
wmHyh8wByI1wn6S3RRRCZYHj1lRzpXXCFPISdY6P2XFcIqDz9I7Ji5orNbhHv564
6Olva/zJuTRV8dRialmSSUDwljP9i7+wNGkE9omwZnbIZ2uSd7CyQ5ihm5qfc9ms
IyQzrnZgAKEW+sSeu5bVPSXe24zHHpnG2nM8/ZsF12yHURb4diNHz2lv6ucUyZMf
7Og5IsYgH7HBvTQJBtk649cLnxDnc6ejv8tQlImQoRtdYK4LTudvOtfuvQXxK6lV
FkA4Ef+H4eCOrlybQu+Fag+mTjWcSt3D13U+V6uaQa901RFIGUtOyH/QP6JZhpLo
4mmCP7bDF9yrH5HGxJPr66cwAdpFSxqxvGCFRPqrqcpa2jJXR5cPMTtLGK0g89IA
MP5QdhwQ0tV+07/yArxyQxked2sBJJzHVxvKbgugQgPeF74pVzR3J45AssWbXxqN
taR/tfGDuZr4LCjnil2ovuXGJlvoFCv6t5GxlhzSvW+kPkIHtBNnX7pIoQ5mX4Dl
8TLfFzZABgEr1XC2KsdYwtx8XNIgyeF/23aXIgbKoMku0NGJ7zzXH0MrSwEMNUEY
r6+IoxpzaQ9XDPj5HmkT4z24rIDYS3859PpBx2+pFCq81Vwn4OnCR3mfpPW7oDXC
VkuzAuxW0vXmGjPtjM9IA45O/JtAkNeM/Q1QbQjYP69QnUvSeDEqhX/Za8ey9y5o
CUirZUbI8U5SWTcVdYM5yHd64w7KATYlP13/L9rpwRR2kPkJ1Lg3jfVJMgfcCGN9
eXxqK51nzB6Ep9rYwDzzJDDhtEShT4il2rwRtYQy0+o9QvQ3h6fG3jHLvavfbT+D
NV3WsEaV0CBLEcpAR2VQW6rgfuaFBiPYok2f10PV4Gq/St/Z77V7AMk6hI2GLrFS
JlrBnXRhPjQN8fUZ0R8mgoITjFsol6uQ2spUi7a52iqZ4Tj0aepXO31bJGzplhmx
10TDMHVUZ0qwIZ7MXQPV6s2DaGjOWbsInL5gzoZ8O2mm+6Povc75GSCg4qGPgJ7a
7HgJ60IaX1IR6zW4Tj6GF0nrEwGZJVuTGpGIqCc2KB/YOAYlM6ll3lF9flG1vXsI
V0Q1bK+tyUc7iqkpBusTWfX3KNZvKM5yR1zg9vBt4e28vGPN5NUR4322QaxyVgCt
598wtJlJXIhlG3Zu5GX/TW77kKxhZHc+Op7w7ngxYUpxz4byOSbRtYDNB3DcggDf
vxaE9rqut72B44ONQd10HzaH9XWAr0iqpsd3M/Rmxwfv35I9F5/waKRQ3kVHZ0Xb
aEzGRCGRdqOWvwXQvmBTiaY58/T5oZJNLw6voHbJuxiWjymO3A4QfdZCbwtzHOfU
WLOE5M5zJ8vpyXt5jSCF5O2QQC9XluBcpT84lV9b0C8lzvnh7QsR0AxuVMbvZP0y
OrWpsxf7ONBwQDsD4ZQ6+qEiQYOSFNWujvl0H8Lcvqn2ix+6b18xPxIQKg5vkO1n
m5hM2DbcMX8BlKLzzWnUJtbmWbXq+YPqSV7ft/Al25DttdZWcOekW/6oDJLnwpts
TPZJAjWNuLgI9yBv3klUX1M5CRH0sbxy+Tz1CGI+eY8aASFOMLiUq6jRMi5brVVp
nAavs5Y57KDk0nyR96vrR6B4xEBSeY2Wjvykrbltmganm5Ar+3hr2amzXLIKKzZT
slzLXcA6AFAcW6FiUMZNC9SgOeNlIUfRCBgGEY23wEa+9WG7fr2ZmYbH2w0l7sf9
VFHmZsTmlykg+YMUAFEnFPWWP3nBRWFtsXYesLaXCEWsd4Z3MZ8x0KIQIFVYnkem
ZiTXPA/7V6xHMKTLN/TXBwaXVFifSWMmtUPuewlk0lyem3yE+VgfCimKU6nvxUjd
RD5OI5OubIMQxzTW4WBlTkiv9/SNlZ3tgVJqSsYHso7KcKf5Ll/GXL/ZLOSUrFun
s2ODz7gCuTDJPpnPX54YFgV4ROcC/Vf2Sxp8A/i53dyhHB6nIssy0XABK/A03ne/
emv+LMwXQRNz4+ZTD93OURu4UXP2H0OKFIIEoE8Ad1Y0GwLI1wDoVok2vgYYIDXO
J5HZMimRp5Jw/2WnXTLZ42QD1PTE7AHfC+Fp0nVmNvxrGiswGzaWShqsjuzPz7vL
o40O85ZxjngEVVlIY0WejzP66rpRhJc/9h8DxsrWBEIwSEDaz/1EeEPXp6PLSEmD
UV2loX411qyZBKQiKPotU7FxNQpZB4R3MA8Xqiu1WO3NTKtnYhwwAqSszzMIsXaP
SfzH6FVg0qcJh+QIUdYtb8dmdc/xrGyhy2pvRbM4ZJeqUlp4a812ce4LZWwurcoA
l/9I/d6mEM70lJnGkeu8LjbbY/8HU9weP4cUw75F1EWb9OGNzycw+UHF3VA/+rQh
1YkCtKxNrsMS8yRqCMbZnlPU33x0NP0O6CCmaKgVYCBAeuvpJLFk9H3Oyv5Z26r2
V9n4UpjE3KAZpZDB9ed3lcLBzO8bXOnCEmCFxvjRycWLpALkSZw45HpFw3hI5eWn
QMqStDTMxzxqQfy0ijXNS6QQWndrYAyrrinirv1ItfOdLzSzl2AqbrMEAcJwEXTq
hec/n1lYL9wODP40O3mSi4mDs/8/5VRgjeuHzQBBND1nDC+ainsFDcS1nXTsMNkx
irH9tDkPelIwFyvMfnSarlT16MGFV/OQ4vMusR+Hcpe6hn7Krs27WQ8/bwrgpkhw
e2WEzrKNTd/Zw+tB/YrZh6reMI7eYAbIVp90X04X+NoeCoZFjSob8TqqgRT2blUn
n8xLTvzoJGFir2kQH1b6BrbrWdm26kKYSS/KLE9Rn4jfYj5j9GM59K/J/nMqsACs
AKRasCzTX7PehPU5FdFNGLiWy9w79oGbS3TDJWU16TKlnByxCtO0HjJfYbPc4B5v
nzAAnAIZMYbGjyhs3UEGuZEdtqGbKFMGRqS+m+tFXP9d7+3lImec/N184vrqzwzu
a6nqamB64M84W1zTjPfEtRUg5eh/8hWGGw6t3nyQgN8irSF59a6QEcC3c4DIh/4a
rDuH3XMGUjoqfcyTzuqRQmAI/86iEQsEhLpaTHJBFDXPeRCM39IqgkX+5NmTPidw
Jb/zb5HDsKQu9rDG1UkgVeyAS28EL/UhMoG2+guy6dH/NlUH2K5RUIOi6Oc/SPaU
ShcjpsFzTZpRoD6GN6ye5CyqILfCmX4h5fGuUbC1BRSsxgxZk70fr9C7d37Kw6mr
oQt7VmDFM8Cs/1aBaEfisiKyZp1rGg+Cm65+NCYMYbIBHavpDh8U50oHiNYhp36I
KmRKk10L8UmD+Suha+cVHBUxXq+UqC4v6PO2oXUo/URNDSbAU/iWdhlXCa76K3H4
UrUgt6+WrzF0CFoYQDivpa4iBMqXNtvkuLgeeb8qj9JMCT5Fqrj1nVflAvKCgC3e
abqxmcPqPk0DDylW+0L0b/rlhDW8LncpMncCQ1IvFW0+1sRH/oFm73rf5B/Us3H7
Rj18Cj+GSK4ZTeu//Yznj7hJpzNdefha4rEP3ACSN8bgjTTiakGTuQk2GC4gTyLY
ssnIXrD5R7ADFLkOYsJqSR5KgDDv4YYmyZRIm0pw/5L4LfDHfQlUjG64AJ/+L6IO
W46nxNMpCDoO+fgfy3O8RRQnO/jdNKI95Ad7yBHIsJUL9umvYewtWgKh4Fw1nmpu
PaDcViR5VzXkLQYw/hJE3RO4dbN/95mLG5IbDzZiecVpkvoBzQR9RuKRMcirqLFL
WLWAh4c/PqG3/7yyJkvQl0MTQcbk2SL+dqFuvEomic3hh5EyXfeTNWRIkAbZFpaZ
5bkem406fHaJvNo92Fy+Kp3jSsALGLMtIIfoEDTuxEbAaH8RPlKvWmhC1yAbLlC4
pUG70w38SMnPQx/YVd+KsE2jwsrQSPG5gl4lxaj6U0EWjbkmWJAIYKPt0YH17q5d
Is3LzYjy27fjakNrdRZZQi4oflu6azisZEf9LVmK6wKlb5jTM10ccYGw567KE29o
boRdUAdjo17SMvA1jV8lt+Bp5zerlSWUWrXm7DQpMYeCgP7eklpAAHAEiiNj7QfG
pPQ7j2z4uYNDw3bVjY/G4wVcjefmJw/FtLkXuC/nblF/rcKUm2i6I8IMlh/iHAo6
QbCSGS0uz4zqhKySfXR4pfZoJKFqovQ50EZi/ukMbHXde58DHVEA2OCmo1GnmdIC
51rwaDs9iUHUFawqWfVR8qHrLWUOLPWS+nWYOploswTwN6shkILPw91NpkmP+b+M
cJXTYgTSHZI36Nj4cQ7iBbDghyv4p+pV24C/GH7RbZHvuM3Dpr8vTLfFO7mbdZW1
Myw+92JqHl9QJqofISe/nkIj51vCsO7vg+frIvseB9zuwVe3zxEpD3cX9QbwZXoo
Jav1Q0SPKXnWw6iB/AkjdwHQ+XzAJPQiBrG6oTmF8/E0fdPeizdEXgWpz4kKNwzc
4qDAzDNNTssEcGsDt/SkvGLzPf9CGnUR/nVGbbm6Id1cCYxwJBjvBcYwfJHVq3Zo
lbNqnFxU9ftWS65Lz3ETHkk5nMhnzkVTsDfvaG9YYZbG8I9YT5fr/RyD7P0XdNMw
NIiUCstnANMHQFUX735sYOwc93Rkj0PMFdDcVGPE/fg3bcckn+W3q6uSDB1OXkj3
aEdaVwDFiEG461/Jk3RuzQtPhcncCMVdfKz9W6ly5I1G56XDCSM5w8PJfLi1bQn5
TWZlbbpMGgzSLgQL+EtyC3VDqgYoL9vDJkWV93v38yg5oYCHY89GuYQlz3K3K1Nh
Ez03NQoF8l+WyCv88d5WWpiQQ89Z8+byvdxxDpN1Dv/sW6wOdoeDMjA5fWOq7srR
0QHmZ5JdKgU2AKVqAMTdyEdyc90/dIm67MY3Fp3cW37rsvbHpGiDnrwgkApD6KDm
Yc6xg8g2qlDl+7pS1p3xJdAA3MQh33g/EG1223IMOORnmWxF37UfyrCP2juFjxAE
QtouNxh+xXRD3a1E4db8XlHPIdR59sVfkonbRD04MMUz9BXqqtapxw1ZvhwV8h8Q
PWk7F2eUtEIls9rdhnkxnLB0vDwLiV90mDe6+gZMvPUMguJEHlxYDMTPA75y5U0v
u0J3cPqg83okvRu3SigD34oXe24hziz09Qm2GlFGO6kDOkr9pDO4IseSss9qFqwN
azhjnNzNJBXdleTe/YL0/PYGSN/0/QSMnCeh9ZPpRvFcRmYBah7hfzUqIkM95FGo
ImkXfO6imcCVQALBd+bcz3ou74f53S6r6i5+1hMIUGnxMCblThc/lsFDnZhCnV85
00L6D1Hk8aKSHESWkaMVn0hSsSS1eUsfRof0/gX244ZsUsoOgjERRLR63UdsZfu/
NEJwJC25vSpaCHHvzMpF2OoSGHdB+daJ/qArON3s/Y9NSfwLcJYTPsAlJ2Jxz3qH
mulzXCq48oNlm4yCa7yd0EPa90v+YpErioTTySbRNmVxOptbApUCJ3CigjRe80Ow
wt3eCBVPJ8UStgMEfzHJMplLG78oyMCrOBYiZAi0oe3WXz/+MQIyPr2EoCUtAroR
jzCjl5ZagHdPtlRLSqmwspDLbH3x/nXIlubJJqG4c4ZJScRo1M/QHkXZXffC2Mqf
WCSJ8g4zWE0lLxWD5MYVzJtztAitdCKMpMel7UB9Igh2GPH/BzvHS+2CVa3THt+w
eU1dfsxBpSx/gH8cAy17Ne9raVIUoIYA/aTx6W4+itMWDdWhH9wzcbTk3Wuax/AS
KDZ4VwB6kZeo9K9O42XAXkeQ1mxP1yBM+trkjVmlIw4p6tTFma5DE2Rkdda2gwYq
YOnmz/Yuw2fiEpUOTMUcxeANMcmTe0rYIvGZrEC8Y3TP/P7t7oAgSNw733MYZ4xb
0fMPXzc25XPfMyouOUP88h+G6T8PdcEZgvUipknyLZr4sKq+PxHPapubshwwzt1C
AhJaq4d94/B43j8pd4zmkUN6lpe/0xZ9EJD8/2btPrZ1U87xpQ6Sx5KGPEiVu+MC
i1ygVT5rjQDIegv7wVJFVVwUAYhuChA+e2mJ2sI6Zz8b6ENJjm+ARoaIaoGx0pv1
ejGat2/YYhSYCopInhCsZP1U3eat7xJdfhPkulGMJTf3r57h2xo/uatDMW1nZdnJ
OyLtUlMED29Cok+IDVuYpKZOULVcatB1/r42Qn6BWS0pY+ErC9yfZC5We2imKVrm
NTR1dm9FsqRPiBHBg1pMdclGcO94O58skueFLTOOFJc7WL3i1WFQUN6VjgMstkHu
FkXY7uFctFLgQepokWQeu5Vnt6pFE+vJxVrO39ECUmX5JWw9Lvj/74KufozRlwgL
rMnIJ+deb0YFcQU5OWRBz/1Fif4i6kyr1Wj1VpDcbDRiBeyvoSP8iMEsOy6SMWhc
Wap1/DtttubEUAztiL4J81AsXEFe57c0TkMwKcfd9quwOJttA6iZzowQwrIZQpCQ
Rt+2nmHPwoob0ByycrfaO4/ZYxkoszDkNypTB7dHPC8OVo2z9GSgPDfWoQrggPmF
GWW/ZgO6Z2svNIJbuSdZmeuQmmjpuMETB2WljNprAEv1g97bRG3mTKy4KBMP+n+r
me0ldC0ib2vvbN0pRFFvXhZ2iLVdwMmDjJWKUVTDZAkWJXJ+tO/DD5wMDcY5QJH9
BtJJxE3Z6SZ/FFTVqBtXlo9jBMA8xy3clAzyfH534/rym+Iqr71wbnCZiGSKna8r
Egqu++dE5iHyW6H0sCPzS4h6+Zgy0bE4Y2tFHh/6OoaUUipR3imnXcH6RqvOr+E5
+Kpo167aTrbHH2S+H61aPuD1x6u9ylrff4YjODrhgMh//F3Yw7DBRyqd0GjNtas6
qJmRFXZBzXlYUUHfvMSyfas5VWHdmXQus+2Rn8gNua7OHsYoxy3flXNcrd+0jx1P
rL+e+wqyrXZ4arUK5SGT07Mgqoy0tB59jjqmz+GF9WorUvy5bfqSyEgh8TdT9TgD
wsy7K4//473mJ9YWppySA/xhcyz6fe8RgnWJAdVAaGiutz+gTvL+eQJk/5nLoXPr
5oxQcTh4RrhY9eyiyVaa6+HEX6aqlgU3ylRy72Nr1WMnVGRoOU3cK9emAuHRNW6Q
xHkSwlDlXNbD7Pl6aOaxNBU9eSqYehXcvctbS6rbQln0GCN0JHrPkfTJWj+6C1V1
RGJHJJD+qivEiP+ELZYUJvT4BhwNlI7+nLQ2HG7YaIPiZ/QzYoG+M6af+hEqjkQ6
qmwl8q3BTi+Cjn0Vx2QZAZgJNeixL0c6Hj1PfsC5ulyMNbwlUdQv8eymp1+wGS8b
fVCfuhqokDwHEId/w/EedIUF4+te4Hs8Rx1iio0nvC5BiI0CUTiGs24Ezb6y6ctr
EszwuSml4a9M0UE2jfyZKy3MGAhI6Btkvm21uIf0AwTV+Gpibn4hk8rpXgH7Nxnv
qi888/rspczoz10GiMndFlqzrxWpzbuMrZ9qWyqpI2Lx6DbKWiA8hpHFdE6YEXOy
Yp20v2D+WOAHXKHbgGgBZjel9gkNS5KnMlnwBXLpX7l7h/D5r6fvMwyZcdTn/uW9
c0ti7cQ4iuXUh2PeUslFksHUyMxhPE2Z53BE3dElk0fNmWJurrlC0YNqVorKQNk9
K1UYD/HGOOhft3c2EuyaSGXehYGhZkGtRtamE17setLx2UMhSXzSsj0pp4upaSaQ
LyJlybic/+uuIafCgTHGmAdCKzjT2ArpdFtw3TJAXuZHBaQLT88Pmc/zgV+J66zt
4muASH3w7kVxAoON3oJmRBCtxialh5E9mpcTQURAWDy4OpT1k2y+ylK1hquPDGDA
nSsydsm6zeoS3eBA7TUv7Cm+26S1ScWzkuEp9PBJhy00MwtRXLBN5hwdEmCIqcW0
f6wT0p4Ya4TFAa/Ky41QkO5IzyrqJ3O3UUZ/2WdNN9QwN12/KZH0nLAnu4QiAXXB
Y+JCiirt8LYqI/cWrxDs7iBRpiTtCrqC9NaR02FslOUH+bBamy2T3UkxtaSDVYtV
SSs5B6Hopn0hhRoMPVSGv9ELtq+hxIwFNWqs9OF0eeschp8NK/qn8qWZlw5hl57+
fK6sY/9kfK4jjkMeMD2hBYpf4tDmmldFCuJUIcsB+zvSFpIDwDxVt6DE1L+dDXDT
myrQMKCoNJS+CPnG4+eWNqQiMuprjFWHKLGf1K8jnpRIcOVwccE2ziWF+3GDmyFW
MS5c7ag6Kdi0J+eYPzz7XZcX0OpuIwZ1Op6laWSwHY9g4u1htNPjKUUpCdJ1YSUf
6bRtgQ0Npuk6gT1lo4bHrRT6YUYjXdseC9xpi5SiznhUEmGRy4pdRs2OA/XnZJKF
zArx6ISu1kshZGG54BQXM0qTh3Ak27LJ6m/ge9uPf2vnOcYrs9/yYo52UBrfaY6q
OGaP30RuDRE6KB1VR14eEGev9Ho73deAgpUhxY3lglrMtZdRVBSUrrquQmSxRHBq
G4J1NgqEgDnNIl8qgvW/KxEyMXcWNU2Gnga8x/LR5Gf5NmyLNrt8Mv7YSboYiXNB
ckRq8lbBUcw2qqlUcjcuCbqs7RLvo9DKcCpE0k7y3z30NDOvtOeggGGAy9ZpRKQn
V+p7SKB5rmGm6aV511d+mVAyrWoDS2Tb0hhl8Fb6g1A2LUhQT9XLDk8FGKbf6AoF
AZkobHJGV9zfEP/o3KdBdu9o1bVrBdqheQif646etigiNI+yYrj5m38KpSDDPOWo
P/8Dk4pM5GHIe1DPJUhXNqvvuOP9PBn4eTXCwcHzu9iZUO6QzPjEulqh22QbgVp/
BOm+UrI+HreqRq3VdCN+HZaklxskTqA15/U/0cIj6shgMgTe6OtQ20noB2RxNaJx
nb+8N8uoOdXFCZdGq+GB8p+EWbrKuJtnNfkBhKCYt/4M8yEImAf7AX+V55hlkv9b
iIPmInTYZhwXCCU7c4A7MVpm6ScK+v6Iroz//nfdoSv1klPYA3iv9w8UxYmB7zhr
U7P+Di64OTivLR07EckgyYrDCcu2XgeQbrmolFrfHnnzOPh/XXXWqZKUSqunR+7H
lssRrP079yS37UgMbDkxLcptXYDFhM2i6Xu3iPWBfQeNdF1bHAP6Gl+YiWH1V4x7
tdS0M4bh1v5cjZeBe5Vhl0b5qhPcmuL8R+P6pDrAv6mKvWhX7n5VNCViT9S8I6Dx
XDMiAxZaH2zhQcJMksNN6+J8H2bITBoU1slQx8DDs3dE5Q6fuXb8HDmeunBB7Q6R
KEP/scV5UpKD+RNywN2DoCfBLvCJkEk1OtwNRXMM5kg63KKcW8u/jCz6eC8Dc8ib
hv3S6xOua1VHRqB0mON9plAun0wCn6nTz/z/ei1viT/LhDLx3s5uo5xUYnKi4AAG
b+li+Ho2o0q0aKRqaoobT5eNJr7uY8mDvMVDbYutmTCDa3CCyeh8W12TP6ADDHEc
kgZYBHVlxoUhn9+28D8ACX0dg8anDxrNzKQx+P11xKpENnbtWO1PiCfxxLHqysNu
uLr5L2YmCITGNoBWB2IcMovphSZpS0Q6DjBcpNghqaSsYGzCBRdmVpN4U0wsENsP
eNeF1SPMFdxOwl09D9hkOQuSDk3YoVXoqkx/fpIgrQWwIvnnM1qT35XHHbIBkQ6i
uOjZmtedvB7/svxPeaHCbiEdg1NqYY9+NPWI6BC8cskpZF3WQ3Mn9MV5IctpsWbh
oiTAGGO6khFaHG04UtHmuBN/Diu+JitHuA8JMqreBCU2Y3/oekbdVh2v3c8lOoux
WVRlYxWczTXk+l2A1JqoQMGrMrE5ZZXfMzj5MQRS3ud/gP//lgg2RaYlzc5m/fni
wfKxwktIFcE+MoBca4X9h0PhjtAHvePjW4hlvm4nn1vNJyhHek5IdBAXXUBoGnO5
aFywgWnjm9dp99DGPFddbNAq/nT10D1uT3Rck1P4LEcmSjR4+q4LStLlQQv8jSok
Hph+8r0lAZMqC5tIj3GBsmNu6/e6JJmJzxJd3aiOxeZKeYS7FKQIImPscr9oQl3g
A3M3Z4HlzMz+dLECBk0mOVpvLp0hBd/lgYfu4mEzzT5Qr+aXSbVHj7JnUBMAw9db
yxUK9eoHXUqU+Jux1rkoE+btvmO5wr5UkYIFNd2PhQ4FoalKgqGdGGk/3ehfBlC9
3wNBBtimDVz8oCUb6eYmDyqTQrRckT9pXZ/eJRMZ3nCpavV4WUCBSFazDPqhBpB0
kqirdo3BjfJWJpJIrB8XkoY+3z27sxz7HuCZyRbUCxNsR3F4VTi4o+5+E/vLM7l7
2aQwNtyH7/cUtCt6ZPGXucwD4W8ay8izkSKSENLcDPa0KpD2qKBD1AD9SpKT7EZg
NfPsUlRHn7iUJsnVxGobwOgyXPS+WH6wOytIzqBiwJn1OuK7/B8ZX/GIvmuP2qih
JZz46PS9dodKpddlbAdy7TCGqQgQ6bLjgGCuuvR+9OKAiO6zajFxv9wzbZPGla7Y
VXKugA1imsaIWMywFa66whrqrROLTGizd+lLYW/51OuIbU6g1tJPDa/O0LJVp5kd
4FWQKtdX2UpJEqqBJWE2nv962IxjEq+ZbWxvHr7VW6O+DqJ8d3/HeXvLS7mbJQsp
qrKnreHgWnF3w4mWlp+jfhd2HA/dpDpMMqSIEhXTJA0HrvE0hBIM9g/Owg0cyQB6
47W/wnevYg71/203P+oyyeyugXjJ/NGvrhSjOY4GaLOoZqfpc3/TEOTGKHv9VnfT
QlX91pAzyO5FviYwRzV0Lu7yLQzSdqohho815s6ylRqLAveTMhZoT8bku9y4+FWt
ZYtHGtwUeSueDeHbslctWiCx9bDK2dumACWRPS9CZZarmcHRa5mFnaiDDExZjWzS
zjFf8FSeO/OuwBaYYdYSFFqeG+Zc83lWxKQOHbCGFKPelm7cmUbvYRRguZnCzvj5
PRS0llthNUcsL5IAp2yEViIC+9qY2co0MM5gLv5uhF1oYI9HlZps6iTprrXZLae6
PGDruH0runYNx8vidvg5dxPVYDegJIyjHYgNE6IFGBxW+oWdFogGd8Q1wlp/oKuZ
Q76kE+Lz/MuWF6FhrntGIfztiaXcfMJanBq5GBkf+qEbbL8yL3L72d3CkeGjqA7F
jglJ96v4/zM1qE+XzORWiW064HPNYSRmmtcMSPv6LGxt44CFCKfFQBj978VB8mZA
nsEkLI237gsOjzFuO6J3/tLcb/Bl87LteZsLiHo+e21qcs9QfxaFeAaVPdMCAlhi
dg8aoF2lgkg8BAolxNglwMS1HIwkNiZLMZ8K7dJZaqLXfNTZ33OlaGBwOl0VIYn1
RhWzf8QEcuZJEfTMaPS0ANC4N7es3KQ5nbt6SZke927yvdcOYKnUrIIkDKG0w1p7
9tlOE6XDR26a0/b1NhT25NXAtBTBHCyEXyRu/bD/2Qxr5+riGaoML6i/NapVXpfz
9/nYhH47zj7tAAjtI/Ip1XFCrbc9XJE0NU70c8ZRDXYHt0kCMo8rFgQb3JPwvl9v
b5Ve3akZqQ1Yc5ncE4wnOLe3rBdEYYQ8EFMi2f++sAMJsw5WMkJhG3N/++anrwOQ
UIR5lFif9qAiiy+5OQqpN5p6pEx0vomDyRAb8/YH9b3wU0GO7ZDfeuQ9WPzoEE3e
UUnU9SdJnYAzDOzOD4BOHJbNEI8ouRflaAG68a9P5XHGQ176iG2s+jTEypLolPGo
lbX8ODUwH/d9GPU6aHRJx/AHJyR8pkqQZc3NlLijz5dtL13EXmF6D/n36M+7oMlm
cCYX9W7ZHQ7LmHwPF0CtpJmtiFzqGmNRLRIFbNkr5mau6WnhR9BP8eh6v5eElsvY
sUv5eFzl8Np2T1v71gZux5HNQmvisL11gRUpItv7qL7tcjsLHi48mKN0+oEPVnCZ
yWj/N8PNsydQbMvQ1yYrE7bvyXh/ufbNRxbchwRW4rIGaPQgtHcW5xE6kW5nGLy0
T4zNZvHkEegFzDkAVQ/c+1RJL13JYDR/wDO8x45Dp9yWgid5LCiNC8i14G/4io3+
AMpKICTUBpwwg51zzgrl+NR3H3pfuWgfATUaYDZYFesY2h2pw+A5RUOuPe5FpPBa
YpvKfbsrg4SHcOvOBTaD4lGBWkgPzd82PE0aPhfSccuaVJ++1L5WUFcgX97Bc2Rf
6lAj5uFIFjGeBJio3XO7l32jOT6PUaLvU2B0Ye8aNvvB9HTrBeXTDlWRrGvZjoik
N9oKZomAa1MJf/BGjqL0rl0TLFjUbamc4XdlIhblDo+iQ5XVl/fusBdMCHtGaDz1
hmNhDgnfuIDdRupbcQDX5E6rMkv6x9IxLzMo9r76UkbH5SaSOL1wXZq+sguVoQLi
EU9po4N8H1FgXLFJkyR5JZaAIeE1ApfSqtn49saAjV9WSH+CxHkKEk2UegdpxUr7
bcyUmYDVkpsC/chALEiS6Gl0tdsse1X8V2p88U3zZIfiHGD0Nfoy0ead6XpCIRC6
kmYE8/N032Jh0O3iZiRiOmPyYE1FLlAYjywvVgZgz1REp+7gzR7/tq303oUaX6rM
q0R5cJwblbNoYPljizauGNPCbQ8NbBTWTLBfbfpmN2rkqbAT2z2S+yS3x06YWzXI
4UVsv0nNDopEHQvYAtY9VKUhKXZGcgceZrW3w1lICRh0O3KCTAlfKzCI2AWhM+L1
yMpouDPJHl9T9duNVyilK4hCQWiLIvbMOcNww2VfK4gpRzbRHdTGbWq450dwg9Vo
9PdydMv+FC8r3BK8O5m6zZJO9mfAgu0nEO72xs27BfLsItwK9PbUK0m7wBCpNyKG
UaGIDvRACwVbxJYZudeh+aU4GlJ8MH1V25cC7N/mxv73x9vMw82BOTSJ0vfJdoIt
bEmKX9UpAOPwJ5RGYoym6KcZs6kg4KyAGPOerO8dopoGqnh2ez8Co0GR/ZA7bLNr
w4IODQIw6JcvYpVNlcc3FZRc37UsCLaiNKwtsN395eD109mDbEnJeYKYUOkLp7BN
6x2h62jw8dclIJVvhH/HH26l8i8ARCo8wlQyEtdeTU8IecdtI0gr+Dql9yRolvSx
oN/cHRoHOtZsB/DAQcx9NDAdXqBCTQRs4j8r6GqibU6NyVxlmseg45mHp5dV9rB9
GRDpV4EIsKLi1ZGq4ked/Ba5u5PsPlpdpjRXkMK2BUan1EWvs+HnhAQOXJPHE+r9
i/oXo0c+TJ1m0JzV8yyo/qJpds3cmYhJkpw5r3Y0tD9VEZNVfsGWEqouak/kS4I4
W47OBa13GyDpzsnWzHqG6PsAFFmkPcBaHUxAN1KTUx7LzSX2LjOgtin+meeuFI0P
y2KBqRr2kQvQlDyd9YYSxHkKdBsLIkhpo8L/a3AMgtROacrhub2+j+aYj+jRZIfU
Yq6HKBeCwsoaechendFFQN2xiCGL5VWCa2Phvy+MISfrwW/GMz7+wJku3S4y/qWb
ivqfFXTS5zOtDzxxiSBFz3aNm4jqXvsFCy0wmHnkXwvyqfSaUZlx5Ltc+P4mcZ7l
iYgcDNJ9agBefzoqNpCWI6jr0+Djg8k0qG5Ag/vKv9qm2gxtmmUexpLrU8X7giT2
ZcMFu1PjvUxtS63PcAPnJRUuJXDx5h2EoZiateqbVpp5CqnIk42OKcHcBQ0zs2fP
THjVNAMV2W1N0dG+LBqTOsVYvghFA61Mfc652sI7hr4rp7Db45tqXBHX6/UB0AkV
q4l1nScjCGF0pc0wwaQFt9eoC/+KRxRYLegJmUKzkYfYhD3MUO6Gf91PnK4Fw78A
78a+1hEZ781ptU+rNqVHzKT+mYhXtVuktpYl7dSTgMm1/VgRMmqx1XmJKXgyJU3j
QBrrOJ9CH0Zxa3oC654Jvyr1pgpTrts0HLEpRdnNen8b2Aicd5OO7mYJ1hSoheyF
EH+s98FpCZyWTj0rv0FU5Upb/9fp7m9GS9zKP0pA5oA6Vnek60WvqPo6f9DQVqih
JSqatLmeBIa/0fxLvXHxWFmNC/fqNS68LlZ+mooWb5UhjSGQdCR/6N6KUNHIzoJI
KQ/pk+NTvV2fpDZPbrEongiBgBO9EfaMDiKTH1A68wrANJUsP1mhpkFTFeErFL0+
mRm2CdkNy1noFMNsGhnluSxhiU8mDsBy/K0u1T6bKZoEng8IGE7/yZLDokZ+Ai6Z
HJ4Sd3BsG0k47L0SLxl9ROxetPH/cP1KCTrW9Kjuh9Y0OxduuZ2JzSmryC8+mv8+
7ipY+RkQOF/oFX5htQ/0A/BprcUNSy2KMXZwnYGuOb5w5BBJfI6BIk9oOO5fEC3B
dAJ4w1ED70sWhJG8YO8TAy2jmrTo44iv67gFqjT0oWxhEId5QSneJ7ja39N5atuA
PDvvUX8qizkb9vbsuJXZlQawBLbDYTEPxkStp0i2KoXNEpt4QpN1i8JZwgN7kAuX
nQdl1DC2kDvPp69jSfncnVFg1ddhvOGRSHx1VPRF7X//TuPjmA9IKTBYJNnxm8qV
FVJvh5K6gTE/PAlZqGZANdcQ/I01U/Jlv8WN57TaLqhX+24uSMJnxr21EGPGANAq
MZaTiuMvQlVsEmPspiE2JB+2lNVtvGa7HMrRt8dMnIJCUnSXbmd4ZUNEr85BN5+8
srNgt/VRpirta4sXLiBM1pklObe2V33biXAiXiw4Yl9LsdCceAzEcI3aUMuLDmRG
Hu2B62QFcVC+mxps8KRWBtHooiqjeofMXS9CQMhzTvStEPcOdQqTfIticxHzaikm
eiLyKI7rPv66tfVEOD1I8yO5/hDVDQAp4kDaC6vsRlKwA4p3KgQTJnxlVrJelHiL
Mssl8tkt3wN/oamf+pM8as9Y+kp7HSTSYJAMtyF2K30FmUviASEmYZvhSvYJkJ3v
ukohOfpNlInDDu9mdjj4jt2MCKVA4z94o3KZDTK+eFjvHub7m4L3HOSY09Ge+WQd
S4ydWH/TUlSx61RniHloTnkUWY8rUOqwEm89PXZuUkMG9uXyWzFyrV8eBi6KYS7H
Btzv9NN8tdNCoGf9EgEx0mfyKe9GX+oO7dRsRmSZadCVrEM1EudMUoIko77fEwym
pUG0PIcLfU6piBYiYp/4x2qyx4YnUtkzjMWojyJ6DycCdTQv1QHKgABZTgEcpUIb
9kYT+hlCgudVmVXoC/LFehssgxWlxRsysUOQtS/JPt5GGwKTSuGuxe9V0wLrNr3v
FEhvIRyXFDYtZcH0KGbBAyddL4Fsdndwj4HKX/HevIOuFJwJBAWB5/ZrWkS1TY2e
ZB+7fbkV6O6cCcpL2/ByZcb/1cANZqbdlXQw91y0aRWZAzN1z+vHRADN0WDD2u0V
zB2T9LZVDBG8NoHsrV7TKqNVq221Ll32CPHVgH7J9M50RXfOxXJsuaTGfaoB3hRW
bN/W9W4BLus1DKeKyeajt9TB2aJOVE7m8zXBEr1izXMTzlxUWAQL/SipofIe3J2J
z8l/r7JpP70e9JtknIqET4wwnfsCkv6rj490mbCawB0M1+DhCMKP+JO10DFPu/lN
qZk0dC83l4HJVcqgPU9qzm13dDXQoK7mJMMxZxFt9/e9XjLqxFaZPpZuOLfd8ecX
NjPRwcLNmdKiAqVTvO+4pKx6Cq/VCgv09zW+PPvk+YEpgc0ZBKWeQGe2nLMpi7Un
oJClvx49XNeiCu67SdVn1FuO8mMftn093IrVsA+jCFNHlpIJLozHncLyK4EFFWuZ
ho23/DYSsPd8ec8PexkeVmN+voiU3kAp4+BDumQATYdB8Cz+IC79dVxJMtKz9TQ2
kR6AKt3vIUlIO8UW/wj173R8slNLfvwREAuO//GRbDm4Jq9wPpcPjVSU6dQMr3In
UBR287QHK82ZXtSM6IsiRkqaFWe83YGJWzNIJjqLwfCsau+S8sn//Fc5zunEnICT
u0UqMen96agsoPrt3lmYadxM1QYyJ3LkU3BQSFVeIIS8nGQCYSVebCNJX5RqFq/O
QSmaGANJUdzssiQK1DeaxrUQsfQKMLpxklXPNRowECpJ+4eL+2A9P6heCCiI+sLf
BesUaHTu9G9YiMvrysapYT4/ll6jS6wBoyqphrzLi+yrZCqfP9ibcjXYXJxdUfqx
aN1re2tV3u/ArMBR//VVSIyebeWAbm+bGNfG0AvaIANCTjanLXXg+FSf304a/pV7
/024eXsn/2syfAzr15TdKKWJW3iveit2wbmSPb6wa9kWXlNKypCwklP0o4FX2Amm
WPF36iUjtgJRombXZbKLF8n8Zrt17UWfYdI4Rhja1dZX8e4vfL7OGKIP5CoAZWsT
q4IcBluQMYY/JEFKsH59l2mOGispl/yQDVWQ3xwR3c+nXGUeh4Gh9FE7/B95zzsz
7xugX3lrByhQhUuseANCDZh6lF+KznRBMbnWdP/TA3crhF9EYgYLCvJmQZQiy8vd
4DcdMqFew13c0zYYWF5/dXVLnPFo7XA3VnjQbV1ZOuzIhRF4VUM0qpax1aKh6+UF
3hGVVmXbMJ9pikUL71RcMfeSq2eEBUPVXHuwFdlIkzwC3DI0yY7GILwZa1CFkWQA
SeIXupQY+Hwr3GRTm4pCEks8OlaU98zqGhua5RXUikPXXByVIsGdN3PuHiVFk8NK
bAwGE6vtdqukPYIppmNeYCws74LmoyakJY8s/lsAJ8AkH8k36OvPeqVeV6vArkph
Pq7IHDXSzioIIqLYfET22wnJswFT7t4aRrxZj1QtsmWCn259OSMGpxmyPkuH767z
9aeaYXvAylJf3bP2oodLQbnkvsgpKoeKwRDuHBhWsxAt8iLV3JCXd76gAyZZoE3f
Bran1cmMnd3JMl7TtEgNzA5XRC4wwg/4LbKCU1OAnNTROLUWQKx8FB+bsw477YpH
Z3eZLISk4gmW0cpvDyPXS8zEKpiFwOGBhP1j4gt/kk6jnQNSrHsH5VQGB/VSayym
Ud9z8Hy9cTKp4MpRuI6JtXj4aA+XENwJYQ3nOkPMyn1s9ciotdDPewPpA5XdOlwF
HHh/1SRb29FStcTKaTFWFABuSOP4JsUq9jdQjzrdc2Kek5Bc22/y1Ydop8GNOqyL
HkiFNQHqv+Yv8or0sdIyDRP2gEmNVdN0hoQuYfDwoxYmWPCTcCaQ/s/po9aXNmiJ
K4kCzxxVxws3tlv3udflWyapVWwlhIFAjFn/UkmguFaBAiQ3YykqS2BjbQ8L9Isr
2l4iJ82a7qo+/jJO4WqLTlzJvEeKyqgIkRgVuabS4mCKPKIz8jfvtdIY6vwcr9aU
KS9uE6QuPBuBVp9zpMvLYY9XIzP0NA6DuvwftotfVTZpAl7wto7qeA78+7tAsa07
5l3dz61PzRBCoYSLmtbOF563zEUHufOCyIvWDPjOf0gx2H1oQV2owi4eYCExtZqg
+LDxXA9d8lKqXRnKHJCMMrn2htbszXFlGtn7eK3pG4KEesGdZBPthnPrckitirJp
gb741UfU42aAMHg/HvSwA9M4tCxDPny6PpynMvJTeXABzpxBytP08//goDKm8B/3
WSkLds5LlfWyWci6yJhjJ5UYzOY4gVVQ29CY6Mk9eGRx7jl+fNoRYdXyjTsNmdNq
RpuS7G8jhZomIMXp5J6UBcbFpJwhTmbo3CSGp22HV1Mn+SZzpUuSk9ze51hEwPRQ
JNOxjmQPaCGqfqPXnuNgrD2s55YOpT5LgG/VIgfgSD5uehgpE3UrizaPFWZBvtrG
a2UFvBXPHas5A1n2zuI1+YR88id9rCaXlIejF4vf8ZK5N5+uvKvhT6ep8z2D1lR8
JP/7CtRKEPGAW0VqCmpe3+IZtd9ZauKxs3X4JIJ7z/nIwGXpa8GAJ/9Mur7wIbZG
GGIZNAB69xFnb9ox8wlJZxQzvBzhZyAm5BeEXsEmW1G4CuEBqFIjgEVHybZ+RMCV
CI7vonh0EuCKDt1kg1noH97vN1vbqwwW1DteU7GO66ay2Fl6+cQA2871emRFA8Dr
g5L+TMwx9BDkQQhui3f1KAdF9e1ojLEgxImGFUk1CGGd5W6dH/mEdtIbXBgu6lBo
/u8PAveVnvpLhpeXgxUuadtka+nGn1QUirvWlf3m4r4rTw2R63Ms7nZfBz3JFFg4
DZX8XlnySUM04iYS/bTJpctZDm+E30Mlvt/ChhDzYcTZ2ZtHPpjG4lSRIt61wxRA
X5+QPY+tBKkwJ2rN89GyetKJ6eLj+QqHcB4AB3/rfARzEhwVEunos0/y8he7Z3NY
w1rvzh0gKf3CfA7/239eoB1398+vST+ZqTNrrMMYNoU5xfq3q8saQNnmVFVB7aXI
LYOAESwej/xTmheVSzvn/ONNBW8s7Y6cOu3FTFx9HMvA67yxRda+8ltLhpX1oZ9F
1OD+6Y+1U6CzfoqywWJ8aemuPCzzCco0jkjcKfvl/WR4KIYeFqTqtMNcFDTqXNOL
C0I2Ttpmkfa+iEyFLevu7MfmdSmfVorqnuuBVqkqUZxiqYHaB0GI0F2TXx8Jr1B+
7vze6najs1Ydssze1hLJjqa3yGuN5Z6QL4aK3jYNrg7tgrzIyNNb7R69OWi2leyi
d/7hBlxCn3T8WdBDIi2jLu2HeDF0zPZYnkmaqu6/y/MOeCuhy3kL8SHDoQmV/aoa
U8weRhv0fjU/53wRc0CBi3asTE7uTE+zE4h5whrYlAXAEkQ/HeS1dlKWS7jrDzTb
7e4DnZKVa1/z4RVrLjg/m/QAkuAi8aBICv2rXE9wmKnBkkSh1yoNFh7LHi9X6LCv
APDD33JStmtLcUczJug8HlnD33Y+kgT4tlxmL/RO6YNLUYUpck+R7xLad6UmHoM1
ut07DReP20P3/I0V7woo1hghA1/PdNJvK7f9k3IOzSfvDuwi/MuALsU2bV+LRMt/
nTTz8A8Ia/sRsNfNoLg/H6Mooqbb+eOFo7PCO+yPJN5WozuosdGmvXn0sjEN2m1X
RscGMBcbyCVzKRqCBliAwASFNYSwKyd2vnIssWay8gyW89m/A/oHaFYgarauseby
Gx0JgXEZRD5tADXP2k/4dRy2fMm5Wk4T2GT75O62bciyZJlt1wMTH8EYzp4adpz4
AWAQQNlvWPClxPCp0Cya6FX96yarE9RJ7zyJESgZ68a7eDxriIf36ASGFd/RcowV
KG/yEOGaBdHgd4bGBsy/Ak6WaasWPchEHcx0myzkNVu90K7MnHyxFNq1sE6Qs6nB
TyZh5Y6Ow/fo5Cp5kaBcKbHimgmHoFVJTS/hzXxdMPuCjXosIomUhvGRpxOoJTFC
pNmsEkvY+HUVSucQrYW7gq1x+8TU+ktHe2/Kyso0hMk53IcxFKDX/GyWffBsUowU
wB7pWPxZjIZn4QlGtiq2ypqroQ/8z4ZCGivulqr8p1v7ciFdOLN1nAMXpn2Mu01u
jtivzeIK9oXynyE4efB3XiyQG2oTjZgR6pVg+TRfh/bU1bIOSJX+EJuQyhv3K2Yt
VtQ5vZlbNkTf+ULS34HEuo/U3GbJkCasTPiReU2hy0BGplSQwETg3wyUT38G9iai
9Hnq7kxJ84ScDgRZKVDR8AoxtVKBFB6ASNYxWRVOyzB7bR89ucu6N6zaJDcFMZM9
gBxQCCWv3qlBnSMec04IHAUgoBI0mbJsvXJ1EMZ4ZJ9m9+8bHey6FFuupxzm50Zq
0ukfAAikhnCFTEv41xX19sjeeY9xr7N76KwBpermCPZOAsZ/AVOzqJ3pK/nvsZEz
dakA/6V9/wOIx+RjYhT0prCogYRUhD0JeAqWCHM3KFriHgxgTZkRUkBpleiC1O5u
Sw8KegHejkYUmKbv9hMmmKiU6eiKaAE2pafouexRetch5dJBtGuyHgALqjXR0Vxd
ou/6FylQ8vB3AgC2qEnjteLd+tcpvKNmB/eC3x5CREpn9QPoGhovvDt0WriVVIAk
0ECod5yQ+xsjF/dI2CWryxwu2vgGXOjE/auPQVGnz6smY6Zf/7cbFKHSpYN5dM0Y
nop5CMP64s2tqtKIQPpgdGGrYTynL9cywsNx9TfSFxXzt+Z7d0b6wRb4fAJakqI7
Q4+EUv5t0oMc+ywFRnvDygXof54BuGlS9RIfs5kV/dgh1QCt0SkToyFxbTb34z/B
2NBmkJWACJx7I1zt7oeRZPX1yfVj5LPE94IBsmaBZzi6VZOy5K3H24Snngc5HDlC
uU+Gm6KTNIQSoHQ5Js8u1b9ptaJ2wCQ6JveEvnbqQvWUUGnfkFGXnKu8m6Npdvpx
LquMADh8qehXJGrX+tYXrLi9EZGrbjfsI2u0FmUq24/WttpASg4DTwpI1dDe6q5O
WJsLK+gaR5eEJDJfM5YQzYhV5XV3W8yTuNTuffEJVzxFupjLO+XFGjKAuL/ofvKK
zxjBWCF4Hn/Xujq8vD8eFV1dokE4b09YqoNw2nc84UvddEJyDXgwY1X5oLQ5bwTU
ZKawFfftWbzaATwxOBkY2V+HG69MvnYt8THVbWRZ49RbnpDbNja/0YoW9F2SbTsl
TZNB0UIbc3vk2DcY0SXMxK09qO5NL9KDVx60Uhb6ltq4xgzqSRT2HFXBId73LmxV
KXkG55ieHJ1Hv6oUkBC28a0Ttl5IQrOpMeaaZF/8zKseT+aT4HNDJ8G1JlxST+j3
O8KcZiGWXXYQLAneF0g0gBL7bqhoHAPUJ30Zv0NKjNJJxPx7Wqv0UELcfSLAaBH0
03wIjAK3XK12gutqCJwz+2/GGRYgfW2jNTZolpcHe6saRFTJRcN4n7SJzUjaWBns
1BAlTExN61WiAMNrR82dI904mGaSP66PP4b19YLbP1axxWo9w02xnmUBZhkxTXqp
Su/CRS2ZeppCLLtXO7spGKCGBY1N+kfwfJfnGfmMjX1rxxdiV+ugbQ68UUoaP2qp
yJyXIkQTwI0xIRi9O+Oe9QZTWK2HKj7eD3rBJkdm+Awq+6ZZu8//a8mawIaXNPOQ
Xnhzgc2mHUrZheplCuNM+NSjOyttWsbyxWlMZcqbBTsIEU3bSJWNHtUSQuzmc816
wBOA2K4OgHWNd61sGDyAXfvrcHTQ2wrMJunlRRf/BqZvGNJyjkVSKyAE4H08oyaK
7i0Ify9j6lvC5kTY6oNXtHDYbspIbnboHAtNxcKhrrukDSFnqC3+/eYmpSjAOHbm
SHETnPAXLGaaLeQnYmAyb+swHG6rVB9Tcc+54XI00G5g2pH7nTBj9k8nFu89JER9
iUT0IOk9a4jJwA/ou9TaQl/3R7JCgB/yOPuLylmnoLMTE97haT2PFDp3/LL3yZ12
5R3Qc+lD8QomvHE38Vuso4qeswyDcFCdwLOCLZGxvAJb3JwZES2UjTAAd35gD0Il
vhT93HWaL0OX9EEO0N/i95OErxoBKu23bdzDQmbCxg6dqXKefOmBk0m/1Uo+IcXS
2aZyuy2S74oKaCLw4Muflba4+7u7qsLXEADMc0w/D6lYpIkXAFbbYjocojgAetTD
adTlI+zIofznpAdtSHUck1kbWtc7K1RKWaQeVnpbchX/va2+O6+NsI6qaMyzZN8+
cU+argiOGTbTsPznn4M8STTcpcJNd62v8ga6wuDV+rGX5hwu59bJXxQ1xqYxtTHb
b5fkK37m68R+oeXjugIZNj1QjD2d7okfF1a9i4/XlOlt/sG0BWk9OD+s5kpGNT4J
9WHT1JdWrES/zXDtdFAcgpu8r12b46QeWhrA0p9Vkm3uGHch/KXitC87Va0p/H+x
xBad+SncCN9i+dcefAW3p0MJ9JRgwOrwdg/LuoPyHAZxBkgBEsRJMbvO9ylYhPMf
1NIiopmFSn2kDtQ07iDVgHqfV9+Gl+rkB5BWVsMfntAWhq787/J4BDTD1qOHrCAn
ps1uFRSTgaJ4X7N0ln/qSYDBkV1noSX9FKOKSki95z5Pr8COTx1gQe7KRNa2KE5q
wRk3fRfpn+xpfuYPj/qP0ZUKpEIkOib7ckvBUXP1PTYwOfezNZcrqxEz5WZhUBMe
gqPGOiKIle09mvsxHc6QnXfXGaO7q4ViMqF2F8EeVdUpDIyrM8H4l+HqGd/HMDFe
tdpz/BP50Sc07QUGbxmDAzbpKujUqJ0NL/X9CLXB2pKu7AouWoZWHua1smNUJiOh
Qdmdw2Lgxj9bI1k1qFiWs6Ah5+Pc1iZysJZBR1VN/eBuSYn03z/D/Ku52pWcvofZ
ObSV/NkRtfP8g7hLWXquCf/OxjLLuH9i73PS0RHAe89KfyCC4/AR6ck7DujzFBqN
0KWKkPZ7Sm5sYzZEAIqu263J2VElEGwAkyftC2lNAGc0qKGCNW9x2uqL3cY9fEUL
1XnJXIc7PrkN9z6w3gllAf2E9uB98imf9c5+SfZZ+DdvaAZSk74vCG6QiqWFWAKF
5sHiO8HC1cATpAiEF82AiwMKotYjAjIc6BI+ACFUtNhHtP9NcMWXIJnzvWNuGANj
1H5AkPYPWdAqHeOeqVXvK3GeTlxB891L/5yqDC3ecyMvHnOZvYc8JE6BpB0RBNpE
KvBsPIhMFjoGpVdH9Us57b9rxQ5VrZYXxp0U9o7RSf0MmsHwsDDxqeopwW7zFrhy
B9HbevOJ/Atds5JiEE5y82Uh7CAmSTTvCHDsRYgIyjoK9YV8/WPayj/W4JjoBk7R
VJStnjmscyNOtu7h3XHkTuaPLVpUj/d7NRZ3li3MxtTuo7iluBXG9vyXuVD4Jydy
lGBUyQ4RYuNIzv0XYpbQHd/dj4I1UH/AwrrzAyP/HgeUB4JRy7YKBoMBqxo90rik
Q9LKEHvIBI8tGLJXHB7aj0U8MxEH6z6oOG+S1Kthr4Vp2nEHnQBo+gStSc66DCM3
RcdwDZHfHoSCXj33mqvGfQsTJEiNXCygmAiTLwdULGWodQm7SGhZ9x8UGCGadId5
ff3to/TArOxcKeTbenlZU/VvB0bAtKaHDK/dkC5cOGaGkFGCGrKFJO51CA+zd/hm
aA0rJVzZsPqUbzid45wA2iw78HNtl2R4C/eGQlPzE7R9so0D7aWUW3smmlPofMm6
oczal1UonIZ/TevD5NluDfoZ3oG5IM/Bev7IYEdW197bNSFZCENJ2ZVlZD3fLXeC
mdcMhM8wqcGklhrh+9WI7GxEUjRcy9H6MOCvkuuD47wY0XMjviaWLIJnZ8TJ4Hyc
hmRcmfECEgDPLUM79m9HA8x8P8C2uVb00NX4WZ9sTcBCz2unOJcEcsQ/TcB8UWZc
bnFsiSiE5rrOMy2didZGZ09qI5y1oVRQhfCBjKhoonvVn/lWA2O+Bx+ySQPDOU/3
yHfLufWZZd3zK7vhgWXhSP7gcD42sfaWtUzrWt6qtWczYxLNCLnBovKc2/g70DJ7
StBdLLfttjw9YoP8K5hhvdZwfBVXZnmNk6bBTm14S07jOF24kCKzetComoPcu9ea
+oWkJtfgg1JDImURYMGOcJ8rB3xiGyikrYWTyhMkIM75IPfctA9tHpx/mrl+eyBe
3t8H2Rzeq5PRc930a8DK4mpbinpISWDuRbBsULFHqrmB88m9jGE1WlWw9vZVAfCe
4GWNwgm+9yg3NNgNP4MS+eMx3rCh6hjHGxw2gOpwypxbaakUgoFFXrq/g4FKhl2x
J+Xd0kRFaBRHTLwvOajbdJ/XfdkDxjuE69A00odOPGEm2+TEo47Ek9FmpBoi8QCm
iN3Rus31DWXL/WrQOQ0dz50RNWldgm0UQT7eLBTz8Lh2L91UccscO1m9ScrpNWZN
ajgUa+wm5Z/p4qqonHOjhCicA6+rNJ01vXgWyeJuAF0sU+W1TEf0ZhlPqGFwTOPm
rUOI+72t2OL4Ed9VF3pZethiwhMUv1KXPrRAPF+y6mWMNJcfbhQ4qxy8d//G+lSB
JkODxoEKMeSkPV3OvI5jHVwj5A+lZXS6X0Y1PIR1GP6MeF3c3RscsoUY6DWCcyyh
BGGcWrbw0DcFa8dyPT5K2CXAhihMipcfNdIARDvTjMNcbwRD/G2Je0Z4QR3YUyYm
ebAXCvIvZ9evZCv681zxIXSsh0xmW2OFv6CvDMiyQmv3GxDwWv9Do9R4RsbiS70Q
Pngr9mIHN0MrA4GHSvTyPZ5bf3FvNMpnNzwpfB6eIiAkJzNY8t49XrF7CaQOzQ2Q
ENZrih/MaLZTjAbXUlnVPgkjoJamXLtbCEyH2pXwWVh+z1PQwA80+kWVZwfNV17J
1ojLMtZwflbPXymvUmQSlwrxBMOSjm6mDcV4xd2KEFN14aaOCHnLMyf3UISSiv2+
3qSoH7jxceKM19eSsjHqa+YTtypxlnPkmRRmKDJ6MA0KeiJyP9ZnjtIzRt7RaXF2
NTXW+buSwc/K3AcjdxyO7u3XIWo/pCc21SIsyyT1R1m+DL/zVgpmR1lWCACU/2b/
RM/1uxTFFW7avT9e4zqZ0FpBdYJ+R3WdgmZGabtumosOEg/2+2xI9GuayOjpwccO
zBqg1RHkgqukuIgDzj0EqYJ0qJsteYP8Y5RieUa9EXTYWBUyaOSdRcbyGYPyvXjW
LvpP6IITyWz92NJJpONGeRX4n368V2qFllwMIwsaSZtj8sdKluMXfqUhBK+SUxRr
iBsQUp8Wn1dy7/PBjWabMLwmoP6WUETpjcRqajslFfTHluv11Rjqd9hG23yT3iGx
GODuqlFCQp9/fY7sRpc/6bCEJQaIKIsqcU/g4MOLmXqRhJcpJptCd1W4W+86Eeqi
Mn4j8WLdb+v2o2LN5Hsaa5jx29xm5IjyyyL5GHTmb/u+WvPJRQaFMz4h49AP6cRP
TAhmjXzZTkyt9uEOm7TMW6PnO1H/Qw8XtHPmOHGrsUt4XdDL25eLy8Fq7/sy8iHd
TzgwDSa82X7KLjBOk9qGWi5272eK8f3XYhcI9U0QNI2/TEd3ulTYUF31BcUoQp2w
Sq/9q4ktd9sl58YNjv8lIMWA4TdpEG3WH5PZKOyDqwQmDdVHpxsGE5q3GA/Ne+4C
AE+2uVgxLuX4QnRQs6OMkSKFzdsiK1mRHDSTNJgitCsv+yG7bmPLQ/TnHNmE8AVm
EAVa1FcCJrkUvmrlFFujIO7kSKWmvSEbo0BtMbgNGCLtsM2QCSjnrc5Cx0I+UM5k
FOpAzoDMpizEl9vXoJSVceKi/YJ8zGffgISdjH9Dc98M5P0JoK5stScsKv+CpH6A
J4larDKLLAdj743AS5Ac6esExI3m/6eNa/K49uqlHs/ZzBY1ozRaIEW3IKdf6YBm
X9R8nfwaQbeOAxWDpjMd+RszhHz5YOGBiXgeyCIWX1ux6q8hNZ/ZLGNyVJa8PDxh
sO1XDM7DnybXanMACgI35bmeJ/Evzha1xkIhnxSonngrP1R03gpiSm0igGhInK0K
0hmNfhenFi+Td/XuusJko/TtP677FrFu4l4Yyg18a1ube3YinUeHzmE5Qt7xcwox
UwgIwT3Qc1lQjwZ1JcxxvRVC/l5693KD2ffQ9sfvnnsfJcCXBllX2Xvl/y2oGpmf
WOBCH5JgCNts/qzZKdS6Qigew4DjptQQ5FK9pPFCoYjOfpCcPmT7M4pUk8UrkkkA
ocmIql8701ajdatB+srPAIwYL/L/Idd6MEvC9AzijIz0FJP0F8uhaYGE6oQRt2gx
b4qnEBQVMrQSQJQi3dXWevZzTwJrJa2hPI0Zjryj/l4yJAB1HdgjGjqtRa2M2dBR
AVSZLE9QdIkkotFpevZpPr6XMn59Vp/uxNyhMgC/nWP2mDMJl/jbe+BQO16yAlyR
KSeWbWCk/fjcPPTMU9AWHANGTjskSKf6Se9UDN/Ng0LyUlJzFrPPeAGgTpmSn0ff
DIWX7DJRHnVsMeu7aQQmsCHzWw6PCiHpa01SSBLxu+mNSjrSSwyrs9auG08KhA7p
7xKz9egjN29/nJk3jfICzrvvRiFXYC1tokIeZu4hK1tB0ZFnNgG2wgWatmaWkDiD
dUCYYn/hicFY+ABk8lE1eJGrFt/s841XuPEjxG9QoyqvWDokwdwYAtIx7MuoU0zQ
l0jbNDa5tN2PtXxUs+v1hVU2D+j90BPXR0R1JNtkx9o/aPJwlkK/E1hOZ3WcPZ0h
d5S46Qwo7zlSPLLOouGBvy89Ia72S7Voj+Zmq5ISSPk/9yN3kLdvzLoDmwDQIIpl
v27S1IXRVEFSnFf4higwB9J4gd21SwY0Y8MHOHR9s5OqB7hwoFLGOKr7P+8oyBEl
IdraHSgE1w0FdXyW8SskA2tuD8lGgV8BjNfv5hPGiaBlRBGaHOpVnrcKJ4p2mGCj
fCxQfKND24/XfWsUyDzRyTf8eoM7SPaDunmk4s+UTvfD6UnixBruYmM3VdnBLYLz
sLrMg7uXy2hS5krKouhbcW72Ydr5qHSL93MZ74FLgn2HKVmcPQycaqmSgghnQjf9
dxQb72NozDx9LXmEic6V0FmfYkY17OZbvBWvCeOVPYvirt5tAc/CBKJ23VZziMub
HGxWD+gtAlR1d9gmtb/7qwIIGugtqavPRt3XyBe4EwCK0x/R7V2+DrEsK7/XCQsz
/r8FvnkMr53/hsrz5qO0uKuq6jZa+XlCwqTJgeZaOK7arW6l85vRREeScpEWYx4H
aud+FbqFZ4zZobv00HhRTDUbnhTYvY5SU+4g+Qx6EyRDC6YaNn51hcVXZHhYKVgU
8Xa0IPPw4KApfpLP6jPXVpS4d4JDYbOPuk99OU6AXEO9zFrtFkw05CT6Y+CDeSHU
Ju4OKEdNjbWjlczyceZLwS0r7wzrl5eRXQonhiHOaBqrloyrtSAymjIBuTG5+Hc2
aI1a44YCADrL+uSdNTehWx8TS4XrMdGrUsmMi2WezCMaXvwkrIpwO8p0NTie2D5o
6amgjJmuiQcPjzvysV3RJPWsYJZA5uJYA1xmpx+0PNb3BfftlvzHPHbCOYHm233r
sUc2BZ7YO1g1pVvH4ldonXzZMb8uAqEUq8VvD65bcMXHJn38CQ464ElX5Jyi9gxT
rbAFb0ImuT3ofedq/FiH6VJKqp7jRjvReZwemdGYvpT3Ya69JElexXHP8QyK5/RJ
KkQ/fUpYCAKi3BSLUq4oHjBrsRrtuUSsB4M88E8vfZUAiLT1JJrYIuk2yYbr2abH
/Gt/V7DAWNVlSrbJHQInshk+a+rtUKfkqVZLot5xGnKpnOVfcY6/mi7ZyFL/j42s
CXUFCpA9k4Z/bdtoVGT9XI1sTlMPdVaXSptecuzlvjq9NnmGA/cEByslXXF92jJI
wgpdc8jl8ZIP+1G+NxOaT1ck2WrY5BwnZ9Mp2fnxA/HDF6pF3UEzeiTr8OdVbB5X
7jJ+3eZ/XKFwmxlTXDE/5E9Tllh867PTJYOtBtINMmUCSsw1IaqC17HUVa2veU9u
b7CtyUiPNvjoklEnvev9Pvvtt+ZhJauj87m5jaTkIAKyVVbEfyVn83+euQidFyON
pcghU7piC/OQRnZiG4gLoFwP69RojOld1Ud6g4udCoRuLqi+Im73TGd7PUEKO/vx
vLtd9WyZAzE2TbMms0rLIhK9k++agV/mC2oINrFPzR45545ml2HXCuKTim2MM9WH
X5TbIiYK9TkUU2PQTEW0zJyMa4ZL/SSWiaTg/AbB/ZeEN3p+x0FPZoW4+Yf/Oh+E
XbNKUiS3dc67XsSSOXNUmzMZerOySfOHJxOhnXS8exsZqOkUZ9+Cyx3ALafZFTxI
YUPLA6DvD79+cNzXYUT24G73mRf2yTWBBvMh4eWSGrfnYmbiENcExMcyG/1YKNPQ
W7KC+zRHh3t7zi2bamgMVyMHI3PREbNiXYzpc3ho6OeG/0OYFAgLTZmSwtOVoNsU
xddCKKnZ/CZyV6KlqTxKrXi1nqUxsAQv8oa6J5ks1wr++vj8/Qipt/J0WtwfQl1v
IOWDy+Ojrh4VSg/SQVfu8FkHD9sxU4ZVF2FmZV46XVuowYOJnQ+IMlH+SpVpKc6P
O8kKO791/Vl7vYjJyuntFnyBXkVJeWn8WfOLceY8csujn4fAmyOfOAE+5BJl/pAp
XFDwDMuxouT9Zapje6kwduDeTLgmppWLJiq0BZf71GsUC6m1esBrzo/UsAonAGmk
jsSxGndIW3jdvNbPvS4SGOv7NLyjSUEYsqPih3JAnYbjwKzaZQIGKfN9W/RtXH4i
g+2BHlM1kZYUyYl8G1gygbKmFZeAraUZIuN3hVA4CbmyMtOtj4BgdOsoSlMOScdY
yMX00s1337wL8pWzZx+PHhJUprVkzcQ37Do4upSEVMVaONQj9WU1QheLG8s7l+RM
CfUmCJoWI1RKz3PJDeI4zb+9fA8JxzWaBaXXnSehQFwlvQ8FQd6DbUee3FsBzTHi
nRZg+uu5oZuwet8XRAdVX2BVv7T2ZabRtUCFyp/3KtIjdWueMlm/HSpgj9K4ehZB
Tj0G4ZXpfUN8O4EvHaScaFrsTzSaGUOR8ANabOzqdun752o+jCeuzbavE3yDFLTs
t9lyj7h7gal9I9PY43GrkzDUJhrarGto3vPIrR9kRM+0UO487AlrsyPLsrkVHZYx
CObiVB62XvcoO4/wjv5cvpdkmVxf73Fby5SVSWyGJ1WQiWoUQtpGcs+AzQNYP0g4
ZbqrGwwhH6+SgfUPVIhvzBosm+B+tw47bT3I8dLxd3EueFkaocNcoo2dDJgzrqFp
hukmsV+bHt9Vs5vxd5bHK/zm7wueeYv2f30C9cBRhZ2Mcu1mR44Gr3+nVoWcHjy5
JGCqBqnx1hX6kWEenptlUUogem9sf5LBckzkPBP0OUMcQGS6IjEjl9XvONiGLgP/
4KFC0CtaLjcKSJbFMa/bmPqTNZVeopOHSVR4b6C9T5icEOMpvOJsbI8vw0pL9uNI
I6aRHkicvsVCjNOotf7iWbza2CFSLJAKGXcobC6WU8AYd2oQDJIQwOCW5KFA81pg
Ib3O5UjTDrq2tFmoJV08TPFNiMxMq8BTsQFZ2JzXj4arByKqMe8WWH9SMkPTf0pm
3WkjgI2WPJA81KZokfIYN1UffI5qdQqFhDan/CVHuapBbl9wYAJw4R1Htg3MNM0p
/p0WS88bnx8vJW0nbVdQ+Lnjl4zuv5pXUcz3TVRWHL6kbTvrrseEDtF+A7/cT8gP
DrC9X6fQDmsjfW5/UM7678Ulz80c8xTH8but+vrN1leAtEx7W6uqLChGDdfX1C20
dR0iGtITugLUs5h/WPBaQYYZTugbEI+eGAIxM1O7CaHyQOP1twnbCnsJyXS+rCbH
khH/LCX9IlXnaNiYSA4X6g/3eCIZ9a/JKIzyPwvJFvU5JPQc15KTY/YmAfMoOimp
Mmn9EGulvH6Me/TR9Eo8VrgOQwVHfNXQiDPRRW1UgD4UVCbGEKg3qAAAcMiGhIhR
87tqgSb86th5wGyZ9MPU+V60Lw1ujPIU9OBHuBB10BT9wACXPthsZdcRY91yJSMn
jlvy/YrE5+0hDV9Jl9U+9xkXuHM+uR1+8mc9mN+cCFE6+J2AwL+0CGxovKkaRrsH
Q7fStjFMVvWj0JQzJcBpmHEbWGDgIyvbf6XQM2amgJ3/AT70M/VWY4r4Z8VKkcBq
oYWGLayKCiLW7RlLNfGX8sZv5TsvfeZ8Labv4neaJnn5LL/7nra5LDvBi5M7uDOL
sk7sysXJy759LdPGGv8eLwO87f8MFyfdun+5wrj6O/qAd7Stt2U4cX5lnzeyztte
10vPZBTngQ0LrVr0koE++4uhoG+9w0t25O9EmH+zwF6DPW0/1d2AIz+g0zhPJQ2g
9Rn/1RpmA4HQjf+sDqbnpARkCq2igJQIhdOWpS3eB9uW7GtmROeiu1S4C9wIIjbl
4qavsua+ARU66kmpU2X8pyVIR1hx/8DzsS+fF9DGwl8qLuek6vS9gKZuJ3MpJmWO
E2HawSTo+dpczR0dbJKz8qwbfobPEiPLYsARKT2Ab1Vsx0I2CKM5IfSlJXQ7Wy+9
dF06QbbkMQa/WA1bdUGtw7DLbXnHJ+RQqRYKzIEsjNwFA9kQi7xVrAxf1DEyyyrm
4p/kqzFf//kf/RPhzSyLed+/84xuTtNIjCnJHEVGa1h/jWDs7ziAJqFO4FdxAh4o
o7TX1VckxmkzeHpxInhJlUVIX0ZU1S3PYxA7M7M+/r4K7TmquF4ZVp+1+itAEpPb
osuT1Fk1VS/Sjltw0VniEDXomwScIvb2UK5257kKv3WiaP1fkE/c2GfYjgmCcIw5
suB9komYfmjDdY+8Bp646lJTFKSdtGSp/x+8jU2RsdA8ngLH6Cs6umSEj0uEDAKN
w1TsJQBWt1XKpD3gKmt9g7ZiP0mGcFaOW0A/kBfVdYRkX1rvg+wx3mlwFBclBOms
B9x1Tibd3bTP67XPgnpBqvFgUe18eAF0DBuvYeK7SCK7jX+Nk3ECFGQDYJTV6NWD
T3h0fdra8TecQLaf8fNpWJlr8QLE4tNW37wfjS34XzbX63s1flCFWbqhSKlKPDnJ
YEcomZZQj/4SJ/twoLZsyVf+kIjzdYGcfjadeABwthYmFFHGUhut2k3r2jF9Do3R
xSq6N0RVoy4GQU/a7pHG+SLTsa5AvSZEpfP6iKAsbbJi0qs3VUjT88Rbql34Fsng
OBxBFVm4+SEA7n6x39y7hFnjl+qsuoy1lFdl9mEmJNV7hARun3uHPljpkD9uM2Zj
9wYZa1/0w3qkxFExa1q35pbX8R1ResJfEN3zou9JXr4Sx0vVPIz5ozbX3WyJzbkZ
dnUw5FMukAnIIPkpyXOKVr9kS3e7iho3NJogbsiYGfxWgOmsOlHrNkDyrp7Sl9Xj
zQeR6NAmXZPgpiQecWLhNQKivBtv8oxjVEWGzhGSYQ+Z4umENmYO032VjEfN0K0g
FIGRTkZu9uRrSEh80Gjk2ruaFhQVLg11RYZDwtj+Pfn2ZmGgo9HL+g1V6EX3d0Kt
3gUi/+u2Z4ZTbb+14I3F1o6F9aPQkJLhTiM6qsXJ6BqCJyEAZJja81OegZJopbks
lrMjZbmlgddyZ3mXuuXZ1VHhrANW88/fG8Qua6BUkhO1TW5G7BxctYMmZk4Ue/vD
0wLsFErzbeDVa7lKAT5srMCYMfsAionciLfuAoAcRIVGZ0SycvhB+g41cQeDa4n5
mWGzjvecmeu1RrfDF4S5EMzFhDnaQXlAnU3cYbQXQRBnpwC4h3c2T+k8iddvJfao
oSnD3dbMwLPKm7P93v4IR6m34IlaANbdxpY20u/CqAPuaoI6za6W0o3o0eR/nd39
vihCp16VC1V7huW405qsTjvF44HRFm/JSk2CVVTexoH62XascKcU6STUaZ9RErN5
yr/GpW7/iTWttkN3YoVmcVj5ZFwU/fHxopiPoQ3/B9IAKrdMw+jO1vkuvNF3sRff
Q4XPq38SSD1W9JuEwtGEt7SYtJLib0Hnx+ve855nRL+R5z+grs/Ou08uuCxsXq+b
iHuARyJpPLeBMujAddXJsLmso6ycp79UtQFTmiOb7fxjbJc8Uhe9fGF9IeEcViO9
0OHZyZ5IfLPHVyiJg/0O0Ofgv+XpjYKDSKTHswRkWwXDOhEMMUY1lfB/5N4kv2Oe
lFaGcciAiQPSz7WG99iboAfP51xLvaxLt0J4Zql3QKETryDPwmrzPyttVkiAef9u
I3K7V4fQvFIeuEWN/ULnS8XPV4XZL73Mekjsw7gja5CHxYVolov8VbhUgQHt1ICb
5oJnOQiaay0RsUn7OITNx3e9JNJJj1w9uKhmHGqPRjrYjRfAXnwajSWI1sm4aBO0
X9esLa3OhOx9QNd49ev5WlNkW909dgvuy/f/FeKPTJOwaKzPBTN6Z3m89iIQrIQ2
nerIMqY5TzWu3SYZS6bDG50JSr5Sz6Wmjsp8et+wh0iI0ZXub7OpH1D+SBgyVA1r
fJ/xKeHJVyCgPFxzmmDhoA7cdJlq3Vtg8ZhpxtJ3aZbhuoN4ZI/6d/G9XEHO5Mwg
OKi+NM5UVwb04fjium7yuxmkeWLWvhNudSKIFu42k8GtB0G0Zro8EA/6kKRr4X0k
ZHZiGMUJRWL5SF1zfC/KUiTCYFzovMzv9J9BoYzO4k/w0SE0dhT37S5Y5NornXMO
PSYnZbgcMiFJqEbjYkYDPvA/G4dI7M2humu1IkDDxZXRoAW4AmEXLXC/SYSuZgWA
aPQCxP0MsjTrpBMrdF3NRXYV+UjaLjgQEb3BLSkHzsmtUcICAead6j8VzfkIO9IR
FmrzXwMfg7Wlret6K6JwFuXqMzWwixikhGZEKGbz2i6xYr5ZZ9aaUyK5c2X/cr6Q
9SakVhI+gUgkn57N4Hx7cKQXe4HfxR3WaDE5GouqhLNjagen6hsV3ichKyZX+nZe
dX3VHd1tH78+47xjv4ffx66eGpMxbenTfsWXuqiEeG41eAxoaOsYUPrHAXl8C3d6
DFT+fMhRY8vF9UzTRdjYj9rEbuXhjXY3+OpizcX8zRrRan5OUdTqQa9MMnwsy7pZ
Gad7gAc8t23xeoi4YfjPYDhhzjPsQEy4j3qUEvfLD9jjCFaZOUy8+3/KoLorALcu
4reXoMvNoXxrIMN/lpeqro+wrNxJfFczpxQt0qEmA82rvKLwW6/Ngt8awtaFw9/Q
A190hWtlzQFEXNTvvbLenfu6WTZ5OozcOF4cp231iNf51gJWcwxYkLhirS+bh4NY
KjxBtGQ/si+miu7P8gKjJWfT8RS2kDv8kx1TWDK+ITPs9ttqpIYb6N5tJvUxOTPV
CegIq+KG77rU+OAAYYIByxmHccrlj95egNyEQ0Def43kiSsi80peKdXsObTbFdSi
otdwjakqdaBERurcZ102enBfnAdgUquBOHYbwbEm645JCeDJBxttzDbZ4KQbgDHn
AwPWnK4UbgBsqt+yp3FtZG8AWncjwqv/QvkKbfxGA17HQqvDo2ebTtADQvBdCxtb
ay6EZbbds14+uFVeTG7utXxDyvczBpBZcQHxMZEaBvw2WHvy7g/wGx4dAj9Z3eRB
qTMVo+zvEQzdeocYTZrD1qKr4q4Mb9Rm+36UoW6FShpeo2Qy90N85Tvp/MNr+epp
3TNMztJdxiW5zV6pmdjHpO+IJQTuam8iT7WU5VRovZfU81Hsh+TfVrJiWnwVZLOY
3Jo7bG8T/BOLs9HhtCdeKsCZC4K0WHofoeEmbdFKywilqeJ2xWT6Hm6JBqOPv/LN
Haf/ubrr9kzVFsB8Gdpfcj7DZUtutE2S7u1n34ECDEigAsC9+ju/rnTyLvINNBvX
05akgQInNmJ6/gZfEuy3ziVlWVhinCy1xFh3TmikFCPurUVpONYnPki5Ijz/omyu
4xM3s6dGM0o6najNEYo1jOmnuLIQxmqNAuMFI2mzSqV0v1OhwE+DiuSbN/yRcwdy
BiSoYFczb10iAoXrvolJuziGa2++oucZmLwTH6TxFD/nkBEcUM0NcRCR85SKxZ4w

//pragma protect end_data_block
//pragma protect digest_block
KZrOUENh7wAfRmxpfF++bUuriIU=
//pragma protect end_digest_block
//pragma protect end_protected
