//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DWY33Z8XfbRUmg1750cEO/vl3J3loosxztFcjFYqh9e0lF1lpONbFkDNFIOyS8qa
TNJoUs4T5gqt9IU7VS8xywgLgLGbGujQZ3mdeArdFmV1rsNKgjLwvooy9nCycWb+
NvTi8fxnxYd0S70mHY0cKQecz+0cyCjcvJ8ieBbeJ7njrTqVIw82mg==
//pragma protect end_key_block
//pragma protect digest_block
FnVQvlMzOMt39kF7wlFkrzDzkc0=
//pragma protect end_digest_block
//pragma protect data_block
T7A2tliSltjygATfCi5U/DGpcy1fZ/7Asi867CcDdGxW1vVEMxA7oLRBpL4/u8oQ
7b8n81kzSUI+KFqlvIz78Fzk3zAXt6UwnEDA2ez3F5zZ/Ev0Oj4eND8dwKFBwqCv
PVOSClGRcMvEhECzy639nZDCeaHe+iZtKUDFEI1HpkFRzY/zHzFzKDXz2xlKGwpl
QPRO2VOI/P9zalzlnRTPaYMj3iuqnOgtbOQqk4E75x4WqGOvvZm6LkpUOv4WEIwy
C0+GvvyVdn5oxj62Bw04eocQoiYbqZeFYy+ZQgaSJKOi8apxEVe9R7zGkc2NM/jW
zViUQzx84EG7JaWwDQvjKHbyEtcPUrm9Wvlk36N+BpFkQp54Fzvx7M7M/qqJ7Ewg
zZQrseJZY799qEphR/3CN+91wtEKbXaNejwqNFbnZOO6vDRnDPuajRXuhbg9dC6N
PVh7LffjOzomKwBFx+3QRN9q6xu9jmh5his0/4uH25tJYpz0x5aTlpVFiNfJdnXK
2QO62DPDOmjkVi/X/l/JDY4wh1senpop17YEUuivvKM44DIeWrX4GXgJucUtsVD6
JKzmODMX8HR0gSjekdYn4+V6F2gsb/mulQSTQd8uKpeAV+67PPxWVJQIuEKDrAaf
q/LgpKd3O4HunDLwBcKfn7EM9fTvRX++Amix3JtgGq0m3DlD6+C3d8T6HvnYorhu
CySdMP6qZdmf78itQmTkTCMvW5HzBtnS+cNYvcM4CrmrNQcGox73tgTirDW80jqr
+iXh/npCjdRm81jvbPLpAY5w+IZ6MaEk5UCsN9AZLfgvAmJXClsqG6ia3/DchdeL
UYoWX8AymyPUV8BWaD56H2hGL6e1MQiamzx++Klpkt0ugK0OmydWx6IdKQNQkKNS
uruIz/owQj+SpLtHzfl8tK6hwWmzIZof/rNi3kRQNEL2AivpY+RP8QzQJ5fMHG9Y
g49ojzVnRZnpeJgDz2ykQxy+cLFLvPTGsRHdzhIn7RFRj7Er3rauvJzz3z2gYjqN
XkOqwhgBeByvELc0HVMnMffiu7UD3kHgqJQZT2tlLjncz+D/s9bo8vd8cggA8V68
GXlDLapFGLJ1GwZcyuh8n8JqlrUt3PjK4BS/cOJQ4jmWPT9PEv26gt0TZwNaDxna
fK3Mwu/IZ9Joq+w2ivqSl2YP2t4Uv/3gwpWgUGjvnFx341NqrCQyDPRotuyJVagx
j3UewQ3wjZ3Qxd3dDPolZ45Mz7coDAnN/xtQ5likQRhs+8Mr2hU4MWsSZe/lW+27
0FXJj0D30gIe5NQ4urpOP0x1CZelUXkW3L96Uj1I/gZdnNdCbFZ9zVnnn43JWR0i
3fqRL2NPDnHztl8uOy6YayZWppashHZ0nNmBi9gSizWdu1q6qKRfmfu28COHwJFV
3jXYQh4IPDGM6bbm054b7pjchs0ltU4PV6aSvtS+SFh99k0tj2HMRfqODMvRaZJS
UTW7RdPzCOI649cakQZep9Ofk6kqZ6mHya60WpMsV/H1NhSaNt7flyuLta2YNQPL
gzYvsLYabePUZNvhXijwC3wmyIvKVcq2ZevxGh4dHrB3NVeNv2PwNsuTOZAHdYm4
IwRCv7M3B+JbiuWeaTvol1anQa6WEd3o3i1RQC6PZZWpRO/hAOKdKT7l6jH60vYx
6Y5aQAmpEHoeSvkdM2f1PxMLOPjvuKpnVOCgENhBMXvC1nvr+uevaf1ZPYbQ8D16
O6OwOf2GC9B5CFlE1yGJENMAVRlc8CoDI2jlk9omv441P8eHlVy1glo513iQ1GTn
mb4o5D/tm3CS5uHstMx0aWPkQ2AT6jp+JwMrHWuovRXGMvfmgjlnvK+soX7JzvUO
7i0Jy3AGATxuvs3a/lLBWn1673Q3tvjTsv+q9cUSzFSY5uGBzBRjflqH3a8G8UOv
y/YNBcjsKMK7t8y8ZW4QLGaPBPySSEumIDyYn2N7VSxRz3Fum/SwToSEnd62/3dq
rEFuhHKgo/+kFTAc2XawLP7K9YxzvqnQhLPg2o2y91Bz93HGHLNJKnNR9w5lfiwU
2kzXv6mJ5MmloRGhHhVnnf89kJDuUu8Fe5e7oU/VND58dKY9LU2wPt/yYEe3Behe
nx9tmdfBTwGebwjp7Ede81JS/fU/FfdQnXqQNgMsNbvovrMfip0Z2/9BsG89oBGT
qSN4czDNaHOjdGpzKHPpnNKwIebOnLHHiFgI3fCo/s1d+v6mz54eWjAKI8UlL40w
LzWUCAgVthNiCx254E10dsjBthF2i6Il2qAJKE2ibs78p5EUygDCxkcSwjn+eMOB
rGoXE2smsD2Sa4GOl9axH3P5WhDCqDlAAWePhk0BaOMECb6BlQw4F7dmJx4K4Bnq
cdO4Nv76pz1HQmM/ph2JrzbGiMUYoKHsaTJxOGhn2NTGA1SNEEtSpsWlezevcu7Q
tnwdem9fcsRJH5yOhuQw/ClyNxg5kbTGlf4gMV1yZWgvCHFLZmODIEwiwPMLnnJ3
yHiExY92nlYs6zDf7LJ+u8QZW4hKa8yjIjwn24RANQfMajRihmymVIxHERXMA1+e
lOsJnnLraNHV64QPga1gBXtJFYvZso3iuaRJ5Iflb3B5gioYO8BURGPkJ3XgWEXW
xmWBsdHbEK+5hKlCUzmLeJgP7aOmszRzIOthjbc6s4P1EDjdtHxvaUfl8sQ132kV
UWynvAD8jGqsFpdt/Bq7HdZrswTfwEPIh5JMqHPXmg9FD5Sjs8z+yssDpmAk1lf6
0oB27aVshDW4BiV7qtJw+88Mac2/rode6wjHnmGoiLd0dzvH5GR2mcs3fFcY58uf
tHMdUQaV1wsQ0vVK+Oz7dtY8LJPWqc/02qh/PM/Dcqgj/tpWbswZ1QKRey89iuiL
nahcFYvDn3T+EgPOq8UmVchG5cX8m+WLvajIDQ0G4rDI3O0XaiM6TP3cuktdPWfp
RY7oGCGAR8byoodnJ9tUKEgSayDSxTb/QKHit3QEAE8Ik4VVZ/tjqH3zG7oEn3Fm
1qrUUO3CAq/tm717rxJRoZ+AgJYtUz0zTv+TtdDbm/3GJl3au8D6MDWWaAWvRDhz
aV6TuXqWy/lclHwjy8Xip6binRpjne9CSMVTlEm0sagYqiOL9mq6xBWeDAWYYOwm
HbuL+zJlqNoUDNo7pcJLdq4tdIZuNb/cxNwScVpRjm4bkzkEs7Xl51r+qF2iEKgp
UdUJWRXxcHS4823fwDT8m+cd4LGRZTB1U/6zBCaE3dPW2pOk59hMaILe5Km23TVm
Z0CMRBIr6HsCZTUTifUBC2dJqUUAg+3mVV8D0/YcDPJFrEEEZYkjEWZXvVlFxR4U
ByADcHnmFRipHlT2Uq6NqhnDQK0SBPg6jiuUwUgh7xuCE7jF9jJuGNoUhr8Y7q2/
KSBvdVD+yLnjFE7ietHp8CesOvJ4UcvDw5H2Odw/Ig5BymI04pR9anvx3DpvtcyF
bXCQ9rHNZtAuRC+ztnXqPc9P+0nQjxmt6/LVS7Bq96xotoSWEpxAglp+TGVQ9URM
WacBGvru75gvCxSSdWgQlVPzsDRkm8Npr9mkjvgptkOm+SWPqHT5HJ7olSMJBoxg
J7Voh4/+V8V42gyXeAo+BeWgLP5L/TSQQbCUzjBo4SetGB8ANu63ct8kGej/7ukz
3/dEL1wSNgJtKRss0TM3PfWaE/0v324SD1ZCY8bO3Fc3w3lnDaFPcNXeLB4p+fcA
o0zegulXQY6wqS7GLl9FdeBLyGF2kMB8yz7gU3qIWG5fXG2ZSuzpNDA6WyHIsknO
/p5q/6SLWgzNgXdCwmQMG0Vfn1B+2rrNQZkNXLb17BHWpmqllKG4K2cc+xUwtSgP
nwz7ILkA5V+3x/volB6E24RB5LqD9Q1GXqED6xeC6s4T7HMn/7b5/eDolU9MhqfL
0IeQYasfIVr36Ev/pcRIJXUUZuMvU2VVy0bRjGPJwCxmSDxP7dK18qaCJHs76JSY
zZFVMmwbmiIWN6A3HfDcZ44GDPltfkcR7s2mC3nAnDUHt3Vzj2ZKzvrawL7APdAq
1frYnOV91NpfqvOoRGjxmZgl4ICU33MowPC9J/nn2alvYAYXkAtDQ9oG93djC95G
XZULIm8wCOGSAXSUNqyrkaf0h5SRIhzVrutLeVb2j3z4BX+tQlYk81MF7WpDyMD/
fYqugyCBiOht/puvUa7Phi1EREEVxi3PJwnUa4SzCBuZ6HFlYJv4jDJ3B+RlgG+F
cGfkYypSEycV+bh2l3WcYVRnfmhcyQHCK0V6WaFtXvs=
//pragma protect end_data_block
//pragma protect digest_block
fPPc2tLrfjD5RQjwM/xz+SgWuNU=
//pragma protect end_digest_block
//pragma protect end_protected
