//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
qtEfl27OzXmjs5k1FX7H+yqiHy6i8zNinLh5mevFlDmlIrRY7rPcTQhbWemHSmVo
sqEn/53oidpeNnjHpRxDRLWAP30ftr9gctq09CihAnm7PRJ8Splyxo60JbII/NO5
pNM+LBqIZg6FxmHXOC5qmNZ943AvqseMMACjvlwhiyZW1jZRmSDrUQ==
//pragma protect end_key_block
//pragma protect digest_block
Oxl4riqFOVhwzo9A2wCIkmwubFY=
//pragma protect end_digest_block
//pragma protect data_block
A1Bdr7MC44BmCEO1p/LewU9g++w2trSAJmqNuGenqf+BaxIrhNA5DtR5irZrBwgA
Kc/OgrCmSTQxZlNgaSZsTFjLxeG0LIrUIvaMcdos6ODjeDZzQoWIYb0YdqilnPQa
qirdxpzBFcHZTyUdEZezfvJRYYCaLCIsD40lDF5ZMBz1OTXMKAelqrdPRhIdwWFo
LggCjQkIEqXRvuWInrSsk23eTdqn0qNm741kDFFnxd5diM3IclgHc5VSN4oZwkXC
REd3YD7G0i5iRMrDyBPs0G/jkiuOzjadRg1rnmV1aYwg5cpUW5zdXtoZXDbOGUdx
GTeEidDKuuFCHuO5gLFiTQ==
//pragma protect end_data_block
//pragma protect digest_block
m6HBEdU++oomDCHLnloU/EApBDs=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
pCTLbpENrBneMwvDYMPzLznQ4E0DBroaDNaTKmlk76O1uoBd2ismxFu12XYOXaUN
GzKQdeAd+l4lPS5A4ORITXwCgYKe1t986Qz/GJPuMTZWw9FQKihF2txxdGU4EeLy
965uh5Jz1QisadJaBGSXq7lEmjUyv4BqchvQaVeCyq4wjBBcq50BQg==
//pragma protect end_key_block
//pragma protect digest_block
9z8OIU+NJz0wxMhaispENd0hTX4=
//pragma protect end_digest_block
//pragma protect data_block
GQxKUAP/Hg0tVqeeYHbCIuBEFrWEYQR0xkzA1UJOrVyUfB7sMXc1AZUK1A4uzdEs
DxaUruSv4NMkD6PDSEBNrytAoWCNeqbnKwytq4i4Ln/WV3s1XAk0Pemr0wNq6Wzi
C/JBTwJCKpjKyWzg5Z4p91ZVl9IP+g+9HDLlmMyVvfuEz31M7UaOxMPGnfsj6da8
3O8xV0yo3hG92AjiZPPhybMDoxkprMMFW/1u2sJpFZom20h5JmHbeqg+lfNznirr
Hdy/czCNlGhj+KWLPBGdDRZA7t/4GxYga8TVrIzwyQAwsQBF/M6Lr1esWNjkQMj5
8QC0gr5sGDcm4luGXbdmqA==
//pragma protect end_data_block
//pragma protect digest_block
2nJAuCEx8WEfcU+Mu01WAohs33k=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wVIeolUqnDQ51+O0W2Qyd9IvxdW8mm/+ysjYBSS92wOiyWlC3N0RvAD6wpzvHIOb
51X1ne6VtTPRi2GCVF3kSU/XlHE9wPZlp0CYHlomJWHtVUUZnV/TNBZdDuJiQHfD
wUdU3xq5gWsdWpr6WrZxceX3ozUh1Y+gQreWzddozImjQu/0Y3cgcA==
//pragma protect end_key_block
//pragma protect digest_block
E4CI2Uu2OTN28jcNvueYPh4Cvh4=
//pragma protect end_digest_block
//pragma protect data_block
5d+ligr++FobSv+QXS9xVWLA7qsLYkzER4KSN8j0LobRkwNA+PM0tSEQKoE/BzaO
Bu4AtJ39ywQ4X48zKCupREHhixwk8pX3zcUlac6XHIsez2+V1i3QxSObtptNXhS9
0DyDRmfWBgqaOd0uawdzrYGuMTNLnV4AJpDuBUtU/7NE8JndBN6qEp247gLgHdDJ
OKxR4nOCHJddsnMhxC8HCP9XA4VOroatnh300oMPGTNJD+KBQVDROs1j4uYx81mu
IqGiEw5pk8UQWjK0/fLTtOt7TaFgjDpjwxlJ38W42wOQz7UH1Y8iFshF/JGI2U1z
T1czoFjnHrA8bai3km+jf8I+yQZ9iMX5gvsQXtQLFiEPyHX54l0QxF9wNZTKsWKi
7gmWoOXvGCCCO97RPbzNIWEWDaz4PhwBHWK1eEcLhkbFEyC6mJpgxg8BAQmkRD3c
TWua7j1fBLrLr0lrprYXTx5/Ph3z7fNScvsUsUGsvYd3hZt/t2Jt/Z86r+VQBrXy
nStvurhGlvnGBZKV4uKQHobk4IzMGFM3qTOOQmKXYDwJ3M5iSVyL0oRmKMYXYkPh
1hNENJ/sM4tPd3H4FjF/ya+7JmqrAGJ1uU5idqDcd4xF6bSeTQiEDFGqgWr+fSJX
h9ktSMK7jVVSrqC7hftUrMcAOoK07PFGUVAldxf+VKT0miQI7ijuN/ztDUEHolFO
DqNMELhQ8YmHPz1rmLRzMAZ+fRTvrAAHahZsMVu7NsXjiDh50Ey8p9RMPgge74qi
XvvVa5nWrEs4/I0gMIvjkqsDypmaZUpTN9wC0eNgQqeGi8e/9adpkxleLzNIqZjd
9JBrP2xnopt9EX/NFi7o1kRaBLDlxOTWhkZawUNN0UmFcuxRhJQJ//A8pqMGVegI
/T3/MmueX9HFqL1B7t58Ck90TTCG1hGan4ON1txFycYAh7LNOwi7QFWaNpq0s0dg
Re9ztAFVAZZNkL6p/buZ+3YPexwPhV4Huw3C4PeyimDK7DilMSuykz8yIE1CEcJk
HJkHVBwHse+3UcaF78nMOMQQZAX1F2lCIs61I94BmDDhRd28Aw8o6zBUxg30p8kT
Ou3Xb0hSeeqNMJofKH6+6pEYcN+tB33aHr3lpLq91hwnRaLsdGf/tJpHqgXcZJvn
dgfZjTr+wg/W/cRLPV/O4NeiGYFiA8U/2LOPCj8FUo3SQGeg6trupcV/ZhDHH72v
IYwwIJ69h1Fd9teT9cFsxq54ui/p3mE/yKIX/zNX6XesnwJyjMDpeQROC9rYcSxz
OMTUPVNYe3ASFY9ZuLEsGwkTHr68s/MD7vF62Cv14MWYvVjSYi8WqOZAfgPOkPw7
TIw/K3ssjrC058md7WctOtQtlWjPli1mggiPF4cejO2EVlUubAysbyonl0+5v+Wm
O6E28LV6r8wonJoOHuvEXEnKXrPVrwJVqPIn8lSf54IVjA0HcIH4I/R+3bstCC1D
6PZ+cufB5U11YShFGij22fil4CL3xMu/qfmDfxQ7VYcGMIsGTLQkS7SHrbAx6fS8
J7kcC3xXEE1wvkGKDx0C3UUN9ECqRU8tvqDPWxNGCACEIci6ryYtwyL1E/cym6k6
D9eEypAqm1ewVn9Jlu4rTfG50ss535I/YHdIBtw/+XgmBzI68K4ohT4Nz576datw
4H47yxo1WcyIEa1zXMKT5hgDEM9RE9Nt6tyexgXOuByFHx4laETCysXpGwbzl6ne
3c/YbyBwbiiqJuyxIwcJV4BiW98JmVmlLQPlrGFDCTw5+qVvNLVxUy4YUQXjkjzE
59aZ/+bD7IFW37buKjkqyitMSYQEYeq6rxP2LIY5JWXhxVERBHVbgVOFaBOGnhst
kkAa1wxhHqm5VXKGvre48abvSSVFpYNucVyG0Y4NnbHwtC/RStAe0AG/wLQbJ0tl
Je1zxy8QoeuYbLF2F2xFdRRX3BexxGUkyafc8trXJrxuMKGyDTxYic9HAEwb8uBq
X0PY7ZM+6xsR6Z+pNNPTI92LlDkwbG/9QTri3ZcRZk5f/Kh7QaxNT/O5ZuasbaB8
vlOttn2fiNwaNFdfb/a/XBjszEGZ0uxkhpAB42upnGrEeUv+9Uwx3gE4hrUYYmmm
hYhBQoo+gfj7KW7u6C22U2snIf5MXsp8ftmL9hbgkqm217dJ3oZ049YXJfoMAhIJ
mRMSOeP8Hz21c1XWNxUlZjJgtrcwRpqBytmSu0Ke6KB8Ih33NJQp+cbB8Ier9cTV
THk7oZXTEg7VgxDSZMkLFG/9af1ZyEBv+3fe831DgUv/vouMqa+/1i+/XH2lXXOX
74T+8gfMiPbcGI+dxFwynkL13/4rBuqK/Tjl+dmRE798GMSyTYhd5zhIm/8Uvsz4
RgbSqEmJJAWKJ+Selr8e73xNi4xKnMGje9rVJ+xTbNHnd8x9XD+2LqP63HFQbmLA
IywPYaVGGeLNtLIfvox6KGErCLbl+YiF6YH4zQSkMKNtDCBIowg5UzYodQ7j/hhT
lvyNRnmQ0586NvVmWty8sgH4yAFyYlGviBfUkBZy/1wHogGNLbeeq+hCxInELXRH
LSHUOie4dw5i7W+9K77mhm36MZ+QAfz5VUMKBpVnTzPh2ii/o6v3t1PTt3dZwn0g
IaDLFFxPgRNjZjGRlCCb46exImWg1dVZJZ69MOzCqiRJn+0WHmLqiOKcMb2+9RbU
xiQl9o1RrgZjBVagHmnF+H2teaRivycn6Jl0stvMX5pCUJa8jJls7H/BAdcEVDy2
5YEE4l9iv0+kniFSbxWSbQc+Crr5fD85o5LrATZsEMYfVMks9AZa2UYxZ6DsJNn1
1cww/FtJFC+eoEvq/rsiTfrs/1k+YcEaahyOSxcurgNadBFFxbPpbzuDeToMlFuo
OMcrEmFhoQVStI5dVc4I5Oe0Z43c/RIqLg2OHb6RFbXtzq540gvif13b8paBRsTE
Vfk38Zo3QFC3KTYiOvkorhIq1X2dcBK8EjY27mjgx+E9EotTIAXrbV85x184M5wp
teO4ufwSqXb7sdBCiudBsC3T+ROzZrnEXN2Rc9J6jsIQTuauDYEdtv6kqHk5bK5Z
6I3VnfJaKKGoIJQ/Kl6GE9cJ7Y+ZhmtyoIJFaE1pQ0q5af+E2sFKxIB4yRGqblL/
amaKi1xZ/fIvtemyPIr3M0Zxt/7aDMmOFsrCl+5ocvErZWGZt16LkHq12SGEDEgZ
UDGLlQGod/pItLyEFAj7SoHmyCiVsZCeD481e5hPHw/9+ARuyjmB2G6H/25yU2Ou
i5NwvRHS+r9Y6w4wKa3Ogm4tGEEqz3LT19hRxXBcswTAIR0TnGNV6s4VRGZ6BUxn
8Ity1WncqYmqnm4cFZ3HIuBG7GAe+TI3uWWpIvAHxjh3cxSrOw9vh3MPwh2n0U/J
caARxpJQyBzoSMceMfWFCO53duoaGQR7sAvLpkQavFGGd697OxIwsoCRXY1Ut7PO
L5EKM9blqSkyqMoY7lZ4iI6q90S6foSk04QQa4Lj8ADLNFEDFhMLKPDmJx1/G7+6
8Eyalv1IEGAMNH65iFBlly3nABlt1czyY+lSWA5Kjure4gb1nWyEiqcOEzZ+lQsu
oXLKZskZA9IUn/4OxIJBBP0ltA/CPTEICWY5rIHyEN34olnkN/AdYpuEjr0pvf2+
A2aA/QklddTpUkZSue+OElhcvJfR1A1PJc6ZflvRmdujsj9AHvfrctq3Fr1X3KnI
TRGFn4eSr+SJCnhpRfzrQufzuO1GsMgEQ2ESul+PnA0qDQy2NkLSGMpwU5eD16py
NAGXe+7RFh2bTo4lKzGaeOMB9M24LLuyT4BXYigsFIvoM534XtCBlppXUrUK/wVV
iI9p3vwwvCfoo5vHbpjCQqBT00BMceEh9UODpUa5FjdrWyYpi+t9TIAz46MjzdSm
RBc8cWKaGHxhOQK+WIxjLx+VO/XHavB2vB1PjIKXLdrnrG7iS7vgT5+uqahgaxQx
U0KwbzftN/javVaHQz6z9NbM6fwfrc4TegAeHDmAN5KrdXsyiobnsEX/tGhAIrVR
xsGrlxvLM7yKsiTmntnIMAsI55W822tFqzKf0FU9FrhHalcxL8G374Tw1q5lHESX
kRBWhpy2BNQ8BC1CSDK84KStBVApv2lhh/JZfUpRDK15bceY/fQgCz0TEsMZKTCw
GPeAPf6f0DyCkclv7bzd3aMxTfAdUAvuKcv6ykkQOBNkqVpv6T/00I1dNIyrbG5c
vhidFNLKEwy3pRaORcoiMz8Mq2sG5B5eI8tK8ipI1KcQMCBzRZvGE/8NgGPg6Dyg
67Qd9rorFf/65NbZhm2jucqPUl5uxdqaoRrfEp6FqVfB7bRl4+iIPYF1Y9vKtIKh
TUI0e4UfEQcD78Cj1LC2GmNASFpDSY2AGRlNgVeq/YpE3HyXpW9EVqU1Uu2EhXdp
fKHhJ3qKtlpL9SfpO5VuqmRsCg+ay13WAvbECqgz+0hVdBz7qVNFOxYwmUtbVxXj
vci5Zpvuawea83FN4HmEooV4+reS3sPCrBfu/h2idQXUOCb0XIEvPuF+qiUpNTLG
pZPvxOWWtjS2VEHEX07m/6eq0tefTXskiQN58clX9jXbHD2zVemZU9Gu3ode3VL+
XyFS8V+0UboEFmOq/66H4nPDRG8N8m7PAbenpB2dolHKr/OSzAEJApMqIfBw6scB
kY2pmy99ykT9YjCC2hogCJMfDy2B0GGcvIZ2CZxZ3DWjXJnwh7+3uISxUXTNosgk
0ryldr09Hp57DoxqrQ1JWTaec/xUkiDGdcoPJTygPaDWQeEDA7wH/kC3a+F1+Odc
AiQ9D1tJWgOq7TRVSe6vOsn7nuDt8+lsF18JcDzfiV3D7O6gdz/JvOxCIeWTbPnJ
gn4pLB930cos0JwE2/0Wxie26NWpMETunCgG27wmzwlBTwei/VL0acyvTRl7Vgd8
2D60mbtM2cLseopzwqT//ijPhkz6OCZbn9Rkg22BapGOBOOJY3EAoX3Y+9ZlRC+Q
fFFTVnmCYX/s3NnYDx5grGH8GqpqqJL5mkyKulyfXwSP1ePwvmcsT/J24I+jMmvt
JK0CiB80BR9Vd/4sCr/K9LWbLuXw6QMN+JnE5azZ3V8LWcDBCUVGU7Uk4UvXcZVT
q1Z85AJjUoDZvyWyFMBu1HQlRlu/heFh7fd1owqfhz5nxZrXcTHI3fca2sbCH4/V
DA587StMtrIdD0NSNOTVqziJFbmeQ4Xq1FB0i1EVb4/E1wQMQtLans39pQrvrta/
EwRmJb5RjzpUsU0dFh/28fun2DBtPHm1wBnrki4b7D8NuoN6iKaeC/hklrk98k0M
/NbGU1qFDO4Klc/tONiScFvUna9ZmzWoM790ykYvvdJFC8XzT3CbIeC798a1uvVw
lifB1IpXPiI2CMea8xnh8nfO6dtN5bh0tdmoLjpCFcY2d2L42cfZhoVKjVMmmDrl
ckYLdmVxoaDHrqz97iZuMAH2q+oZ+IaqMhHuF7oXIS/FVTPouzqXyKh90NdhDfuo
NhfNgJcHgvsx26fSxhWsgiUXRCxZ+ywa7+RioKxQ22W1d+zPgl3SVs9lWvAmAzaC
iq5P6PXR3ZoBeX1ByTZ/T3TyePTmq0lanPamrW718PbTSQHbwxkifgwWbIJAz9+P
LyJmna6rf/A8E3J6vkmi4PLMxy1Oc+SRCS74eque/s2fV9lyj8TPoeINsL1Skrwn
HIV8MU1pTXFabUNpcUCjd6dTs0fzCnqoS8264B61U3/AMFURqP8hne7CEk1hNhMz
BGuSdDwzId9MEBeQ0U/6NvALGEsSGZ8fLoJhlZ7w+Pt/01XnNmFfaedMuHJ2uDTs
FqrMkonMcOV3mjAlT43WkgAkSqQHmov5oS/XZgJtlISW1de7R+rjiDyKfK+WVSoi
HLODYKyy3orUAH3FQtwnLq1nltOh8bEG0Hpa5DdMkV1LIO1QjtxX+HDKOV2ZVulr
QUQ06WOp4Cz//baIQx2LHmc/tzIzxpAHtFmGwG3bY5A/W+sF2Wi8+0Cf2rURZ1zd
LZr8s/sahj9EcwmWmPauWDZXc/9fnO21E7ovDASwhzSXlRNdXo98BDrTgsk9xC/v
besW9KLBcwGluZaYeOXgzbZI9urn5+Vpjg65i6OViOAN71jP9/ejaxTQBhWyUu91
ArLkwu6pXZF45HJE+f16+p8+QdZoe4BR211Xh2/OaKjfBt4Kt0Lt8KWaJH+zh581
BZM6jURyAKk873U6qxvqVP+tYf7jkf8767v686Hu8vkFrELPlTyjA0A5Qt4N8mEw
TAzbTERRfHvRzfeoS5acjckg7TF8JGc9axjqnOuLge0akf4qdJY1oWD2w+gy+0WO
WQ4miPdgZwE/Hv0fOtUPacfM/QlYDr2px+eVYyd5XMTQKCf40J0Tp4lHRg7bCaBA
bV94LYPwmV4UAwwjX5hwtVonkGkPyNqIU1rxTJ1fi4EmVUcVcaTyKd1SGZ5IVaNc
UZt3fv1FI8qIuKDN4Sj6z7c7QuYSyMzTdWNW9jcPYuG+Edi/OP3+TH1t1g3UuB0Q
HXrxgqcu0SjUzRR52n1w9/E6yUGP9P6bsIe2uaJc6oARv7gETckkiVoARMxFAMKQ
eVSYXNiVyKUDuS5UPf5kmBImdPbK40bJW4DcQ1GtPo3qxD6FQjMH93bH6L1FUVkq
0bTzG71lMWkzs/yXc1vl0HpH/CW2vpBF5NOCxLT6FYRVwnRTWR+ikBL5kMirmY6+
fRwfjOt9OWZMRpsDxtkkFUklKzaMkICPdm/wcmxwo79Mi91iJ7Q/vhcTQSTYvZvF
LimxV3dSAfPSlq2TvrGEmHvKA4XhKepWVXWYx8+qS7BBR3SYmicemDyNRRZBdLv3
PsQNuNBvUrZs74j6xkwI7S9jO3DPNAL89p59n1XmnIe22lcOW3vgQfV3yqOtDDKO
IGA5RPnMl+ZqumHNiKgMe84YNK56lH1CJ1jAObnCqGkF4fUYPnpKiBqWPNp/9aHf
GmYlrEc0fmGXHTJ/zgjzfFLNis5+uExnq+OSJwXx/sbSJyY9cn5EqkvwPv2lAwFM
xyJ43IiHEzWcVFtuJd9kls7sEcZmOPCpHuZqKRS168GgWemzpCCmmNkVBMRRfHqT
h2QhULjolNMoP0gUihYi8Uy1279bpHMMfZbsW3gDHNwOdJQGp5oWUrnTOTcQPGp8
dW/wOAYYvSJhRRAKO18UP+5pUrmvPSbGgOlU7Gt2+AMuacGnLqQ5+gLdTHFSGDCH
blp3xKzEOVYGfaeBKtYpO6RC42QjmqWQ8xHmdCMUlegz5nyaBkgAJnfozMkAQeos
3FDGE6vVMX4tSCtQaPxoFC9ygQTYW+ys4wBuS500KvxqArzSh8Y2OhQ5NhoRciRO
hHjhKU/xHPyz6WMVT5BNnHe44jCFtASH8KAm2ssmnz2p9WMHOktguM2774GiJqeq
8eV4CYOO8AQMEfhc+XFS9jgOUFodwrq7rLTGP3cvcCpZfgubE9tNIHrz+KPElWpF
ce6mj7p8ffPv8b3xL7UvlF0ljmG7gOtD2JIQVPdESNUP/n+BnqZNGz33MQGFWNrh
3+MhyP7CVCNrLSo1930a1zj+OU/LOw/BFNOlw4MenW4ZBWjsbFJt4dUqcSqsnUlK
ab0SZajK6cn0pDASayJJh6feo99mAtenydEvbDoPe9H8+JNQDzIdSw0PDYLM7nse
35dBvxsj9k7BMsMtYiLL8T9y7kvYmDUHXAYYmOKMez/G3h+xIVKrwzk/OD0KSnYm
chqrQB/ugDHfvpsFJQXRfphKffgSpr5Ex/himuYAs8DyM9VJqT3CCf0RKmvaxd3H
EsN81MD52qwtMPy6ImD/WyP4DbnP2R/INIIJaXU5NaJk60CqLYp9MCSn2M+U3iqu
GFtlvelTdEm16eaUZrDyafACwsP7mMYexT+p+S7wS2Ir+gd/phCmNRnAIvg7qj3L
lPCxdkX3CFiH1Srt+S17XGLTn+eVGZlM6Loh+C34+ElfUF3Idmlz5v4uyiKt4TbM
2dm+G1Orig3BRtS6UnUbnVvmUnAphE1D6P+fgNB3lkMH8+NhehwINGuxiN6cOwlu
Q1iHGiUTm0THekahubKUmMemF/oqy3uh+R58GMFEHs+Ap53Xww9QvNCnzKKzwliJ
1VGb1Z/L3W205OQ9XkCMnts3yxh+gbHfXtSnGPQMVzTbfYvzCf1S/P2EeB1H63GZ
Zq8aHx1VEmH2IvwUVrlckqXwxWYY1q4VBlqbwh7QGJHzYiseIE1ekLxgRbqEjkl4
VyE4K5LgLYmVutdMMVZHxBHwxaxkqUBo62qSXizJ53ENqXrLOR432Pi61TEXgCzv
ild/QRJ7Pc/grZmQVRh0bS7PS78vx7q849MZamgMRwiUZeax5yJklJhCxTXHpw98
ZyKZWwIQColmKhdnjpL5cGNt9PPLQXZE10sScK79DDlYkm6DlhAgqh/rOhF+9U8w
si51GQ8N2/LgWCI5LzN2e86asCb4cv9+TuZZXcNF+UdffSw+VhxpsgUcGSWWsyZ6
y1Zqx8rA1yttMC7CdtshB2oGKPqoiuTWDuC1RHSSlQzwDHF8f/VVBrGt8sGDUWEG
A9cIlTGM2LM5tKkMze33BwLXi58QEDdQxgvk2gCYBeZvC7MaiSD0g41sHQIas2wF
7f/5+CqpxFZKuUsj9S/CKgWwNOV5jSinx/JhK1xvdcIi1Q0fW+lS7CfddtPvV0CT
gnBzjexe1Rcx3Z6I4kdU1xdGKrkZkVVl/yP1gcQ2WyF/Izhl12HNMrayfXf7oGJJ
oZCyf3kTEpBzUxJzRQJUc7ZrOm2RdZfZhcJBlTYV2m9yWogEFqP2BKWyZrcAKzbr
X1NOamVWvSyji5CjUEIB90Meo1uRcFaQVir6X04QiP0Q3FBP/QKypdhjLRveXxq6
h3K3LDN+iLjGxhf3po0B7BQO/tgEIFfk1etL7VkQLDfvlcdkxNMz8q8aGa94E8Vs
wv9gBYrYngz1ndgwOKf4agHgmadNmcBaW4bsgkGbV27qN/7pGpPlpxgR08sYbJy0
EHlRkTSBothReI/F2d69eFoszGxIchiDdlziWMkbCnHAxvs/YFD3EyAkkoWx6Jd6
lHXaOAHuWxBHDiKBD+AAKZxl9qO5AYosYKU6vrCmhSs7zlZlO1MHCDLe94GiDcnj
ZmJpP+gBTpP5D25ZYUmrJrXWDT9DGvL2wRy21Ff5ImUlj7ROGTBPztoHFuC32NAa
1k6PFAaNXBjbEbPaSO7BKZHtDGDO4vPlYRPjmcpKqKQzifOMWI4MavdChPpdEks1
5YsQ9kODVbELu1s/D7WasTX7fjOneuf2MMGAygLUBD5klaQi4k4qf/PyMjllrB7J
orNbBR/HCtgq72WdGKiqeSItOusosHnabBIrCySOr/8ligZ6FKK0W5SLUhoGy/OS
6NR+XFNpf31VgmSNLupAbDLp7VNfWMVWT3N/yLFbMet8tyi0E4uXFIaX49TK0z0+
PyQMb/Pot0GzBr+CuU4fTLvaNg3jVhibvKzSrs93Nf5TK3bh2AedZv6vYQ5P4uag
aszI5BdGXKYd7/aC3CkpY8iviyDZTTKZap8k8STnqlgN9wEY3UrdpSRGvGLRk5NK
PutGeMQYyTvVvs231a12hhYn7qmqKdGz5mV0ZcI27MS0Ux5kHC5AjFAnrEyNLKOU
dmEZLHu0X0gYY2ND5v5LpiGGRhSqRHFsVSUfVCxVzBJsKHIuGHDiAs3g7fKLj9Mp
Kx62u8n7ti8F2R902PqJNrZAgc9GjupcZNSYN71yu3von/pK/iX1xc+CqGVZ0Jju
/5l0c0+XSWLB7DTtdLIA1hQKCF1K65HRm1Dln9QRUqp4Oj9FFkJmiFD5ypM+sKI1
EDaUYck31rBc0tmTfDm1TDveRz0h9RmOfTJL7mZUE5YGGq8ppRo3be1lhEBkClDz
+pV3TgqeIpIFa3wNwV8O4ZZgZBsdaIk4Yz2qsx6qUgXJ5SLXs39CT4hsGHNYq/oa
qwIbLWXirgGDaq2ivbgPQHh65spQ/ophFDYFqDoqdqGgsj9JghtS0wqUVSfoEM9K
4wM5BT0lKHnw4BGGSdlxfF+jXx2e+bEvWFAzWVWNEmHoUdnmQGHk2Y/BByxnHg7t
ir7d1JqR3r4vOdSR7sBq6niessxg8uBD/xfMGAQUiKOtTF6RVMBBfHvG76NHI/uf
1UcI3Wkc+/uVGE34/f+bVV5L+E6ZWoyTBjenfpuHTY5ILrDP+qWQNmUp9jlsmFjt
i5t2y/+XEdHXz+x/eJI1cmc61s5fkIq4FSJ961C3yYMD7Xe4i9uDMNVg66+V/vFk
bosOA5VJNLgTyZRh+v6V6PR6AzuxNys47/lGRmMLMu62zLWxjgwF/Ut2O7fWjrtp
xWvzYUWg5bE7ZbiwNEBz685FlR4sl8JOyfKz2V+Jax4EMgCQvoQ4+4cMqPrkbjLT
PPhkQ2DzKxOivH6XjZiU00eR+7lcuT4A1R71gvKuOJUuS0A9vwCHCOVyFrvSMxX7
fsVORH/9M6+sgjzPOtnRDeaOUsl1eTxPLha50d7Ocpi5/dGEzw2iHxJg+KUxghh1
MGqfGfqpoDE4/pfXurRwKOcO62MHXUottQbyQGasYUV0v+e7Jod+9oPjrrBp9vXT
pAAFlY07JKkBfnqTsfRXVrvBbPBjIqCyknPvIhTomB4Vt63l0Y5tdeIvs36kKbt7
9Di6reDXcMM7Wq8AL37zzYtXCVeXF9jbwMHHgpoDF+9lRRY5NfjO1HpnFwmZvxYe
JXfkFUgFbRfi/MI0pc3qGdJjx6Mo/z9MayB9Ppq6/AhUs7XLaUk/gRfb/UFrjFZn
PGut0zxpptlnzdt2YtgPgp7TmDeYXa1MGz+/5652QlEfDG6i4tYCo+zDe1OsEyiz
ZtslgCHlVthIcqAJ4OMTQopJ0+gLzlxtYhtO36ucYxvjt0XJu2d51AdJ/pFfUFcd
l2azrMzZDvsLlNfxQmSpeh7gEE5KqusbstXBv4/ava/a/zeQBgeQ691sZevDOoOu
921dYhubu/DXCb7bTBYHI48c1Ai+/klzgt5Eumx4HtAzwKSkRKLuQBlyqHf6Yu+A
6T5UPLGvynIg/97ryS4chi4yy3+7eJ3fGQwQcAMIPC2YMlIoGb1ewmOgTKIBZILE
eEy38ma12zlO4x6IBOYxEFzYaaOmH7nvy26vVh4DzHbTpAXdX2RkfxxSwzLfIZ3C
E9YgFVvXLQpHjUjl0fNB4/JYDvBQrLhsyHtuO2sM9DjF2gkfWykuKkU84II6WPQS
Q03a/0gkbL15UZSCWoRdk4NdPzG9NntNv9TtbnpT/eOsV4K3IuN8t3LJiDYnVk62
2FTCcn8DFcaypj08Poyabqzv4XSqLEti6WyGtWTpN/jc7Pl1jJUiROWHDmi5kIre
SwCDM/OjZuyTYorGzKjqUX5v8gipQowMMp4u+HiKvVuhlwSKr5k48JSRMXgPhafw
2sLVFW9ccx9tuRjpp/5k39lKHkEMl3By6YZ/F1+YGxWGfuFiR6wGhSofNLpBZybu
HACCJlxbo6my5CHFNd+eZuwEOmz7i02D0GQJzewt0rvLwVWwEKRJgn/xRvNttTOz
yTU23cCFgGIqEeb0KqtyGLuXzwxIDUGx6+e1EAP8Rp6ZrBxfIOHVImhjjs0U3uFD
1vg1jCS2FuFzeKji7zbsnjtEiQZ432BIeJf0GOhpkwZiiZx06kTDntuHzlsbhm51
FfHDeX4g9bLJiwgPpSHIrJsHlSKxTJmgLoQogTt1nWqvqdycPweXI5n7Mg9vet3+
N3besz3i9Nqw2ekcE+kwdR5VmqS5HUML9SaHvZ9OPddE+qnM+HP59nrX3FsX4lci
yjpq7EyVD1L6wEGfOtyhM+1bcyZoeJ/4xjvPKXWc76YuWBxtkPi46tOChdmv8Bq0
ABDnxmxFcngL/mJ+2F0kXIMWq8M990XoM3U0F9Bb+j9dwPKf1Kfa0OceFzjuJ+rM
qUc3GUPmzS3NolDsGcggsOpPUTIEQrp/U6JB4iG2z9fSZrwIQtG7l+KYs234yaV/
kkUfuAk4VkbuYhMPP5hDS0yfy0E4dlO/akTB8OHYrMCRh1VWG9UaBChYXEYtIFjL
8GFV5rQpWBXTcR7A2AqIEAZnzL3ChrtvQYVCv8O2eg0U7xEA8sVt6EuxBZ+O3HW6
koaHUo4uMr3FLumuA96trlDDXuzTcaqTD6j049zbVfbax5qLgEZz3pli+Rrers0V
tTkPNb+OkAokCni+EscFEen93txd28/5nUcqW1WIkDqo/cyVb2E1xI+eSqmR7v0N
H7K4ENDjL4tskNqNLCXG9TrVQs3En28naE286o0fqFF94wNBzReeu5tHwFCvD5RH
irpEfNUkU1XcOvEI8z9KgHyZ+/jCbBGHAbwoLARxvwwBty6cuXAMkUaDSh+wBQhm
cJ7TLt/qO124qerVOmvr0gxhEeoMh4bV2bHiKfpmWrROU/+gqo6JXLreU+1CPy4v
CqXSBeNYTexBLBrgBROJ7LscLrcJrUMonp75kNoqdblLd3/63FD+o4ko6GGq8hym
hqxzaCkNcQwGTtVG0mSLr8wi1sF7xa+WxAipyW7q5W8p6RN2mqK5wgyqrbnjJLH+
5QU7wnzqGl48Q5cbSUrRfgcOc7fwIXLy6mJHf9KSiDDaUM1/ZSnKJzcQWgSfZ0Ng
DiHgOd4aVYlm5T6ulw3eRVes9t3r1LLvA25eta1SoHqr12tb2LD+htpGHddy5zGQ
dg58EVD2sL1V52qNEJ0nRYB4WTfwRCdZOFoxjbR5lMHDjuoIlY7u+JnWQArpQ9nz
reanWg5ZZ3ddIbh+0Mf0vVHNnWef4Bct1pRadXjVI9xxirz/6guW9mt2Fg0DFr/i
SthNS8c4qs8RNcLWIdG19JQY8NKw2pueK7FurgGGvr/i8gY4ET9JVwF2bFbNAxFV
XoR6odL29rxhSTay9/U8oA2HQXKN3Vr/tkLLkhgeoNrkNK4M8gcFn4MEfb8Q9z4H
Tg1nmnvzfk2gpqgvfMx02YHEswSU66MaTz3RH1JF/iit/wcTvckLnHTsYEnP4I0s
pNotfDachSkGcvD+kTB70uSS9Tles0FU0GPf7uqj/2gVrtQew2igZf8s9woJ+Nmt
UUMajQ859EsTlTSozRiy+trYCxNtypi/mXcN7IJwq37kY8fAB3EA+hIXMWv3m/Nz
PPL0e8tsRTz88o45bTTaW05tIzG8n/6qs6JgyNqXlDOKDPbeI4v45qfqL2sKqTHY
8qvCJsTqE5P6jwPtSjy8kY5Fwb1U8vIPHbX95BQEMhZAINTDQL3hGUxBE0rUPVgd
ESE/PG7y8cLoOlcUOnz7YLfF/Wfy6OdTPkJW+QG4oWsInFW7oQlRyvPaKfQUyTD2
/QQdJUpS+WjE+5y5kC0EKugsg+VOCK3wtiDvs/EeP9hMJAAKLTBGonG94C5smrjK
9bB7cC9WA9oKpfG/1XrO3wYWTPHJiPrpwgXs3dP3aTYU+l/MbsTj25yM3w3POaE0
ODtQ8HqEQfqAZd8oj+XtU6r42/lEyvj0pJwnPDZXlmCVckyaOnoizGirF0Xx1Gfe
Esh+PUNPk0mkkkYC/xbLdb1oQ7DidBSs1Re5d3w3B9VgCGwZql48Z4ajw51St0iK
JuSsn00A1zb5cCdHEcz74ahRdDejyBiPrvFyeWXCo/nQAeIfis9MPBAjfC18ORSP
5RTSL/qELKh+02Z4AwDaNgG6jKqR0a1vhaXh1wPvLh1GlDhvDq9ElMi2YwJH9fD/
YYHkXSaRGmME7H2M8LGnVETaoB2f+VhBc2Wq9WfN2M5DJMXuWNnkKqOqIP86ARIm
HqDaNG+5g4ehN1l4a47uxiNP3B9wlzkYFRC8SiPs9+b47pbbO+l5Ku4CI14ihtTl
Ok8BMpQwBbkay3ZhYCCSfX1HFItTFJTMkOWJJKwyrtZ3VhYCCz2F8EhXpvx8K7Xd
3pkCTrUVWHhohMHyvYMklKQpFI0DgitAJxEjU3mJ04I3agzWqeO3+mUc4e207V6X
+s7R5fVDDLTHwefJWfrL694XzWqebZ9zsmv5Tm6dT0K+inKYQkZkqR+yIcAun0lp
npT0dMNTOYPoeV+R9f8MYodsBsIcrEmV1mFie8Eq1LyVezza6i4NwRrxVadhImEq
VHG6aJ9RqzSVOq63sYOUe+XbG+9WnE77MtEXFCyPKPJm5ByMRWEUOV8hvk62W1Es
mpkDTttuUDtEH0rEVKOh95AWF++ySPtRJDItXAp4an6AqCvdRQuFwAkUTkfmymSP
3zWRVqGueUlclVASgKJyNA92SXv8vGbhV0qkhRY9YHGS6jBzj2AWPUwZfvcoEIQK
wmE9kKNBjQ4xIy61xZqQc2txQGPk4QMJvFGU6NZGLX4KNdOidek0pCoR4l3Y7/yy
NPqFgib8ham/60x4F+PRX+jol/HuC7j8opv54rVhaGvru7H3vxXJemiSk/aqYJx3
iYNmEg7Xtfm9U+jVBBe5Omxs+s4n50/rfenkuQyAJoOafBntvOdOJuU1xPZbuAyR
YOiE1zGKRQqzRlY3MaiQFyRL7tL2SK3zS/+NDN3DiBMMJh0tGBiV6ePNqLzBtRBq
1QVJSHTjLXmmBo8VCJbBt321Ax9KfAAYH3DfrU1FblFDSvD3vaKkpEwPbwiB0J1A
jZRFKtgSRnkbAp5wacGBmD3lCGn212V27w0kri320UZ165FZrKuDXyWd/slvTI7q
k3uh2Wrrt7WXmPjBktqlFGSSPIfbwkCGlp2K9CM1E2omb94ziqhbRit/ExgxuCaI
ATMiGN1IYcAURUBVaHGr2qvaMh+BEKr/IzULwEcUFyIm1CzNAaDhHK1jjm77Rl/7
ifZeZa/rxXfjyIf6qu074OdrzRFeZKqqvRhv2BbMtq+1uQyhMWexDlxEgMjOO0+K
jLYArUCGl1gT2No2Soy4/qmCplFEAJLjZDrRvHsm90O4PYK70cudWpOhF1K6pr7c
fa1lpACszsfIqnTFl5/xPmeVBCaqOINUVhse7vnC+eKHY8EKYtV5cmhNVm4D4FHZ
BW/7L+Ctk1YShRRF6ZvkxUVA/ra8XdwKokxm0FXq6BeAurGYu/R8ouJMblNUqR/z
tsphokLp2w7SbPHQO/GFQ1UXddX1qicRhzKZk/CAFXjr2a3lAB9g9oUHiYJ06ibl
y8DV2awpjUSqQIEXVNdKXUTDtrm7+QLlO9bR7kPJ2zF19eVyqaESAXDuEtZYQFOM
eUBcnm+vjmIxwH8D8QXe8CDi5Iy3kFYPJMPI/W2tUQVTdlURwaO4tKteysSXS3XA
q3dasZIC9wOWINh/VcEkWUCu2xsaTu0Ru4ezU/gVVR4Px5+3YIDVJ+Rcl+GHvBeA
srY4xWEFT9S1rTlugoSQQlj3MqJg+d9Hv7Ey9VbSM4hNiJScswJ9p4aSr8sSaUdX
JCUvhar+W4ZfUiusi30Kdll2wI+2ei+qM7mfVcPP6/MZs6n19IRjqa3Ucef0FofC
+j+rGZzxLjZAGzm2qmTL2PW3srfhNpT6AFQrUGaPO8ECm0WnZZCO4DFNQb04l70b
WwH4RbstqbpYscFG5sPMe1OKtJ4br5kwpB80N683EPCUHem8XLyL1+z5zeDjuvUW
WHG9HllNhTJr23jhSPypCnXPLxuMLG/QviycM369LweufL02k2djPPCj89lIXt5t
v5VAz9idBHBG9c8rHxzlKM9cBMriJE8U/0psnjBCz8l8qaG85sNVpp4Lg4TeVQOe
FMP8pr4LVu2ztqdYvC5f05GBS0/a52GN0TRha9QvM9O042U15Njb1JirtOpuQyGR
Y04GTnZ93zladrAGA9G5GmyvrRO7XIy3OWrcFmeoDbNBCvRWDyL06THl/fxpePdg
pL1pHJjyqIqTNeluXIIga5VLd8OZJIkMileGQkWJtOGFqxe9TB4vwzu8L6FBDugz
V25i+BvZ2wgC/cn7U6mLhqB/9oya39sWpnDuCM+Yj6SdYR/QU701lqS4yCZ3Qky4
++PF6BtcOK2sx/H1FQi3TJs7rN/e7jCN3/Bo08uT73BDZG1tE27tiXU4USf3J1pf
DRuio+I+GOTK/41rQK8aWwrZ/jAYI0B69k4viH+g3lGA32i993LEcfSQh9J9QEiQ
/FOrZlWyaNb/lDfbuk68HiUS2M49rzSIjku28LVRjRzHG3CAHSiK6K0azdUG4C5v
OcVw29VWIMw2FtGphHK7N/MNWaUPfa8JvZ9MfYl7bP+tOeZhCSROKauvbzI7otIB
pUW4GNkPvZP5ROaeulIYo+nJ8gOw2gHPjiydCpFousCpw2TIAiVcWiPoRZmk1dRI
u34RP/UzjNgczqUZV5HmPVS2pU/6JSP0XVhAwQB6rTi3orTweBRQxzZsbOAsdPIk
B+VcieGnROZ/mG3v9iFL6cm33V7CjEkAIJinOwCe5MM2KjIAlU3/f3mkLFkIbHUv
5hbKFDrpxU+p1ILCtEDOp7aXZ1KJilr8bhuJDBrd5eW78IpbFWhIdBLDHohu2jD4
fcthdBWhXmZTHPXFu7b38FLawXKfQokV05GsC1joZZxJKQOxypf36h+F+NQxYTJZ
lhcM++lcJfyPbhZ9WXrHs7bzU5+J5uO6MZVr1OyZgil23nEVV9qUGZLztta4Yxy+
s2fkbbDNHhMXXiwIUgXJzR9+eh7PSwm0tit9hA3pjNC5m27twzCdJmXW1JVUJqqj
yoobOGl562TFH95oDEA/7/FgQhDzdQvDKwsfMHDBeixURcR60RnpVc1wYyIu8ynt
inEDF4VgXnAYIg7k/kZg3CrCdkzlWisTzfjWitd2JKitNm2PEhSU2sx4fOUMdo6I
ARJWzC0Spata2ocSsKeIqvCs1fiftBqkAXCV2IbARw+GeoDqBjtgBgkb62mGS+5T
G4ZXUVKh5JwVIVpnGWbsw7X4czbzMPqg6Li8pe/AS4rXYEvNcQ0bgmFeYbxOHU4i
zqoAZRNH1HbjwRXHUYy/j/eF7dilrretjKNVAZOBrxTiaF1CH7jR8nOjYo1ffSzR
qvwbsJCME6NTz0e+6WHUPOmsfdVjUotd3C6GQaipKIGPu1W6TiQ0wBRckloBgQs0
B5KQOACFxzVub26HrbpOEp5ETEwFMIJuetsarAambaccVHINafXSLRG6AESh9lUX
f538B4dz27OE8VgCSvvWvGA43/cd4JCymRcnqCh2y1BkZp+bFrJH442U6ZmuZITR
wfhhKa/UuubTPRp0xtVoOhmCSFTpzCoI74nktpghUaMvKu7PNtXmLjZW3SaCG+AF
81woASF+VBw9VPo/KAnAjcECnscxrxly7/t+wrErqWDCyLcy0S7D6pwrdnwzm3nQ
k/dURMjXeRyMAdbiV5ITUgjUye2yl10Lxs/Fb6hLfLGp7ONn13V7koqtE+c84T6k
aGkZxLJpeDabFNjXCuyzztw+QkP67pd3CR4A8Ket3Jhic/KFhvdpqbgEh6CW/3+y
l30cSrCpduzF8BIzZXTGZtvlhwTSd+apfa73SuYBFmYe1E3rKSZSLp+ayUhjlFcX
mgEpGJLsLteu/XaGBjIDVGBJ6HfguTV3TsVQH72AkjVgAXTPYx4EJ/an9gQxqxiZ
o86omfT29IsZ9mLb4WoqXdukSDhVOXlU7yPpWJkAg/UHNYFwKgMWaeLSPtB1Gfe7
NZb1K2IVuaQciqcX08h+m42EYiDl3ckofBh+zRS9lU+Kn9yCDhvq2UKi7ZikVKPr
7lH88qX8Kss4Ik0oC1bM0DnrNiJgLmBuW0w9UD/Z97L3SybgugTwMQNRGwFAyKWm
SrHi4HIAUDzSPSnJOgq6Gif2TBgHbR0oznhPCNi2Da6WwAC9/JYOEqhYiNoLDiT/
18ammL5LE7Diq+vXiFN+8tfn2FBi8xXWtL/W/WS8M2oxHO2M7ivILWFJdhrAhHml
tf2G/SfylJSxtzjjybqNncFA4L9jC6sdS45YWWqvs71n1Sg+OAbqztGA5i0OJRFg
JUN8++U5oJrPOR+HueLxdnThoWc8u6hnEJR7rkvyp07QH2qVC0t/yy6ugFvBe0gy
LKiPhjI6Jybfpz0FBx57p/s8n1hmwoT+sT9frgYp2+WTvMVEhwUY8gVS4+x0epvt
Vr0LI8Llu0QkFdPJak2zFdRCEtmimilRb+olSIBW5ZyTrBRGqeV/KYzrTmjpvdBK
zVX3l74ErrS6zI9yv78GcjaKQf17R7cjew6xAOQs3KoRdX5mVSmdMq9W/FvvDiLw
YS0dkXjb1ynPdbDTUVtdDrO26p1jRPhjElT1mXC4xC0lWDf6TZnksZDkt3lz7jFs
lqDHgbbOTG3z7w4ZjGKbly22mxrJ5Vg63zRa2Vw0hvO/Oglhmq+oCp6CvvOVQmOG
6uBiTkJxyigoxUpekwnWZW23MRuE1nlrONMUZPAcddMvxQ4U1bGbr+jkv4868Dbu
c1pCkrcyz9RpjhHv9/V5nNamGvPEWwYnADzbJCQqQfobghlM1IjHfd4S1gSaEs9i
9LeousfS4qjhCkzQ+4NviVI5zgCPYC32fQFsiPhclQh7hmnV76bpyc6YFMGanloX
6yi7idGxuEhM/PYn5Na9hbFGf3h3RAQCZtCMcGmrWp7mHOCAVtvHdW4jFjmsrc2b
dG2suPMWppbp17wsWJmIRYz7aG6VAzSiAzBrQYMSaLa517DSzNOVH9XfpwHLZI/D
jVAspRvdfKqOu5POroBvNwZRpoZnsOXq+RUXd69s55fwvVZQGoIXxFWcEbzCZEia
kW727D4DehLmd8UJxuWYMrBWVv1J8ayu91jeFeOwll8w/RSB0HyNejwzrvBcrKQI
mUYZA2A8D24+Nvn6aDldw0+Od/LXRsksk3B6hKohw9abUEkzK297rRNslez37f2r
p93VlEp4QR2jRZ8kROYqaAM5jjCE1NEOyGcl/xvM4Q/yInp11OXPvqVhuonSONPE
c5WBiE0L1TP2CiGWRKXoXHO18MIIbt5pGk6sgZ1GHcIXrKoZhca7cWv+LG6jfnL7
1MpqHEW3x4V0POWoKu+TbF7uX+6mb79risQO14NucE030VYvem1wk67d3UzTrlPZ
g94Dxbha/Pg5sVg4yKsfA6OD8D1QBWvuhGHcRu3L9mOu6jxLDgpjPMtERkA8WGUn
ebPalB1emcGz8bnEelc1Je/Hju/SZVqKkgd+xjSD8Gmxc4qHI/Lbzq4Ij4Z6aQ4i
Qly/ywD9VhcNVcBtXHwCguqaQAWAiva5SNHHvLihLIX/w0QfFBpD5zIrwBiAz9kH
3Z42qQQHMUHAHlSJEu9+iRr8glxzz/pg4k5CtJOlVY9qpGMortUSFrpBZH9wyMqZ
kQ/gN8lEAemvu9fMc806CVY+NWIXPXyWn4TgwNldWqwELCxk9t6XI/X1zuYyNIrt
iTUkGBmuDLtKB2IlLLdc4tcL4BDwprsDMJ2BFpNW6mAZGPBnr6IcGJS04L3l+VBA
FH1B4EVNkTPnwvvklmdvfufhoE0srvxHVYpcxzmQAoH1hnVmOrsPPhzM4BKhezKO
EGXts3gCYZWT3flMugwVaqFBCsSAfZrJwMthgEz2kEceWg6P81zQS2l66vMCqkN5
O/Ge4YoMS2KIlDn08BeRkgyVZ7WJZv9bj0HFXNJctd1JsxNuVy8ZlwWyksT/xxLj
w59KuOoVrGNHZ3+awJF1OgG+s12YXDfZ4NHh9mIs/PM9qG4hJl0kiKIH8hlYOQ9p
qWGpNGUuoscK52cGuEI1cL7pKMhJ/2vkR54kurINxCPN1NPdxOlBjkQgyEm0LV0p
jDpWDUxQ7AQH9Byiq8ZqFGAULZXXjep/DUhvpksoM2Mhvbm6kKoRhF9o9ct87N9X
KM3d5dKTv90/352PiIB9khdpy/hZkdk7TrhBLXieUTTeXfu4PmxyO+QtmepgIgeN
ZY+iWCFe0K/DtLQQUDegVLequ1o6PQmY51nps245lnhknicY0SY3to/doldyzQ3i
aQ/eUJ4eVYkuGqeE25TdGoRlmSpZ+h5e5WIrsnVQx3/0mv/Zn249kf+9+ronHEHj
Nc6rwfG5FytBHLGCIJ/xGbPL61dilah69VgwqihHBQPEy6z0XPSBdx1jUJQVCACp
8EHFW0u8x1lY4i/m4GGjlT6PVtKkMpRBY2PHF6J8ZVllM3F7AuJmXmsRhn3ZM2qM
aLdlAn8sMRIT/LlFwfFuJzbN0R7Gndm55dcYPEfZqDgFmLMN4GALHt32EolCG5Bp
CBVU5X6lLJAj3vrPNdTb0M605Wqnp/oKd3Z+p8ToH3DHEgWTrvZQz9ZZ/BTRXeKm
R4Fv1bOQ6o1QTd7K6Fv1ui41BPR/4COJ6y+AjkNaHECzGaEFJrChLqnSmB/EDW23
CT2VJUGPJOE12Q2rlob1I0D9WrWKzRkZE18KajWDtYaJCfDawW4379YEru7v2GtG
Wi3AZGW8bFgLAfF8/FJv5vU1hriU1PsilCURyhnfLycBo26ALEPdggaL3zB0TWM7
uAv2+Vg8h8Fk5Ce5ZFm0v4lSa2khfVPPF3Ys4P40yXxwaFaY57tsvqaQj6fce9Px
TUKDyXWDRXTOXtmAwCZ58JpwWEZDqfbvmKX3D1v6nGi2SUSN5Ub8IZs/BTfmK3e/
YZPbh30YsuRCDnHzHbhl5k16D933dau+eAjbTWh+SIYxi4WoOyE++z3msCDEWLhM
U3j5PAhGdVpaCJlhMhXiSQ0S8jgnkMe/QXB/sf797rHa9wKAUjS5QOWpXQXkPPhI
VX8z1Yxa/Jgqx5TFji9F+SCoxglorkDj+neoKjG6dlk+jqDXRHFKmneN130JULj3
NKooz8gHjSeuJDgaQ6BD/hAZ21RagFZHFxwmFnqV+r9qMVdGbxg895GTZr4AKez0
sWbOXONQvfpraP1szat07qumTmfShNtFKOVmHqVp8MsU9cE7KJopn4nqiIZQJ9Kt
Vtj3SM+RmXJN5INoms2/NFsfY1k2wMp0V1E9lPIG+J2IkRTlwCXGALrmwP0gH3Ya
MSpm9/IYmPh0/RkQYYP9tkP3mIczgiOVpZKSNS6SLO3sYjd76F+tpktE8f0TaBIU
/pkOkgoB6rmySXdVJl1hb20dCZZuhCamZQPwspDSeDv1uZ92GiR7OnppTxnF7dtA
R1F5yBwnQX6EzwqaKdFgEeptU4tn8F12R/BVSVb/W81GoGqPBmj4RXmgLgMcOgjN
hpd0TfhhtRDO+Tt4o7Khjd+6z4bzxwMykA2bZ3kA3Jb9+3NnGmwE1e5ymvjotINt
7iBSZ/jm5RlPt+hp5eEV4/o+/Uk6KnFNDZ5/JgXIufdziwey1OQ28KfarQ0gbF31
A3jxNlGbsGvztCqQqENZbwr7cA8cBPu3elLWJuXZnoySmzLYsJA4r5GxSlSMxxix
Ge8UP6nRqt+wUNW5wUJebprn6YgGvYVf9aO+ND6rnxp/iaflPFSjK1VkYli+Qjce
/vQlDpmawiPZQywFF5L3TDwUjo8utkvSL7k0ob6D2m6cCwv+iFjBeYE6uqB+bRqp
sEtj5g6/TP4MJtj/Vg3bcAJ46rBo+QLcDqbgNLamkkhDQCSP41NhILaMGuUpwRWD
5GfK1S9hvDNYutkjEQMBRiBNs0Fv/Qh0iFv1V5Y5GGOtQ6sz6/0hq+IbCJrZjyUe
0/sGP+NYCldczTgT+Odat5WwOEdcG9by8y6prItuqh7teRc7e9E6pWKAQY+TlTHu
EYf7andzSgemJonTla/DMZhju1sHK7tm2eAowkdmjk8ICwR8WxFkeaeKnKmSxfcC
FGLV1xnUHywVHZuPw+i/6AuObiYnu13JcwKcReL034m0KdKJAw73TQ3tIBjx7Wyc
Myj4LSlvEspuiJFZZtOtHRxhBHlSsOoP/jguKF/jn9REIdZLAzQwkk4sWw8qVWt2
OgL3c+nz81HuRDs21BJSslOD48i5P8kiyZ2ZTdCwcmsVpc5lj32JPzk+9/yEKxbU
/KwZJyL2y3tpDl1a7jPbiM8fB1S//Fi3r3QuqjU8jctf7mMO8/NzGkwfB4/SHj6R
ibER7Faet0qPW6HuyPQ1bguyhbhgTVsTtr+8qM9wefe27qP5YRj2UqHROVFJPziG
VmML9M6iufYjfDpfXFeDM8flcuNFKbu2sMKZCdQriC6LQgA0pzEU06VkwkSKKetw
F13Wsaap629GKkq84/bkNkOoJNEgM0lgoyl355S8rYtlcKeKCdMwMJkDZ3c83WwQ
vS5NlPruw2nQQvhFB9Z0kqtyrVpJYO1Lve2fH0zTFiZBQr95C5k3nyEIqlSHyIKx
zM8L350d38d1gcoHWhAenzJGjEIheKyXulYlW9/CRV0aVfPST1m/KXyPZPnRaa/l
HJk3t4VwNz46/oth261kXn7I4onuajCuQraQyloPos6kTcHIhy/S+meejPW3yVqu
T5GttUA5Eps6zy66oMm5UEGcOxZp58FKh7dBsT6fkmcIEsrajTSBNnPYs80OSLo2
5b1T0xEcurVj8THfIxBmJDaMWl0jbkhpGxtGASNFwK5CT4h0cTexnrYMSuCgi6QJ
ooxjDuJRhUC4dbvGVTuj16fTmikM3PjRRuJeajkzRBn6DsR4UE0nXcL1/BMRC1tF
7j8g789VrfShdiCedr5kFMZ0MvDvdhrWnleu+59fxvs52TO1K/9baxNR39xLIlOU
SlFVOEDDUUXlTZvWLRLfpa6HSouFtntGwwLkTjbfXtQADmbsRxndB8d4ebsfvFbt
MIxSSVLduq79YiZLHXoGTL+pKTekjezRZDvFX5Ou+8I/2ZnwAQtJm+E30Qp7SOQD
hSMVLgjcZKs9eFHLac9FLGVwpzRpl9NKr8s+4XKos/rEFZAMN0pu+P6vT70zRj98
Tj1j2HHyiF0IEAwMXU1Mg4OzKzLuHAWepT6yiYbyaej56plMuFkkUaLvWMBfkmTj
7WfP6aViuH2dxmXdH/jhFUq+Zwxe6zwqIh/a3rKCESueMynikFKPoFiVOCK6s7dX
23xcZvYAClWbDncD7jIdnEug37v7JRuGtpnp75ZmFElOXCVnLKRVXqq4emCTGUoX
BSafX1+xv6zx8wszdpEcwesdSP4JZ/lt79oqlHScRuo8Ecz/ReXWZw1pV++sVOKr
+4tyuDijFuYj5EYL37cErsIZ1gEMV3cZLMGDYpzERBZFav9vQ+UjM1CDb/2YKOsg
UyLqe3h8sS3KSS2sIlK646o2UbnfIeClVm7vzDbFPeN6QstHDXtw6/6FrDBUUSgd
Td7YofLkePsdEiX0jFd+hRcPTOMMEz/ag/5jnZ8pfueICs4FzuwBx6chGBnthdTu
BcZ58rUzvaTP7H5UqlhgGj60Pb5Nti8iCCMXgFWmCzfXDZCpB0suhznDNu8Dk/4+
9/W/tBI/9F3k73CGkZYhgMCrwiv+UH06L8+LPRJ2J6SZAVfNoqvTwytQkjaCI2AU
1u8lr1wwMU/ulgYAcTGhxexl4r3AiMuOImJXcN/Mdyeb+QriF6kw89v3vN9yb1mr
Hh56e/ap0F6EVOPvkPHLfsy7pKm5Hz5IYjxkm4boHdblB6+AevBhB+/RIi6agQ8j
xAzxm3MmsqHfd4k6g9aCRl2Fp6rtROO+phz84hNo8r6LQTlYqWOrFduN93/rCTxW
jOWETMQSMKZoXpiXvq5Q/T7otwH0hrmpd1bonn+JBP2QERIg/uwJnYA7GVdEQQmo
3ryI63vz8gd6AgoxXh7HnveR9ny0G5H2LmUpe2RHg3J4a81Q1QtGMLCI3uGRJwBq
KkwulPBG9FlwOOht0qnZTPoN0G+eNKgWGx840j+QuigB0irr6qlFs85ZQxnrY4JX
SVPv2wJTSLpuR/KunXmkPOuqEM6ugj+J6Iljm6yaMObwwpGHcm/zfcEMe2bpoG4L
kwIEy6P+2912IUn589GqFWyFHJNTij29RZCU6lqF0mHzMmDZAI6vE1TwIuiiMMSc
h9O7VYmWu5doRZLorsvOaMG4K7i7gwrFGlnZ71o1ZzW0EI9SyMAmnYDI4svL6iOW
2xy+1Oj4gwejktptoei/QPrF6wL4bch+7zavdA/YScNbDuC1s3cw7MqwutGggnrv
67raZ2Z/B0vRwvIoj9uVEXwJWQEpwVje3ehxe81ySoO6RES7rhm3zKrECK+O3MbR
2S7F3YZFXJlNFyjZHx+L6sKgtqzxeoUatLH2KVa8H6RIUSVVPrrgQSpNIy6WyukM
S0B4xZUIzf+gYSg/6GNc5JFe9ep/iIsp5Bf9kYDffPuEqPSOaF7zWotQ6q6lgzKz
YIkrcUU0NZmhCHpZiKK6NXnXwzYAyeeNIzg+zKd09F+f+hS791DUcE9mmC4z7mc4
mBzR9puu/hHwZ4H0jPo0S43nv7OUwm7ZTWupEcjfctBRVwFBcXsVS0ctV1HPnnj1
LjiDkE5Fd7PQ7l8MbnN1X3+dvsrL05RecKeDWX0fN1ozacsqbckgxk30iAQAQH14
reJMS22Q52mTpRWQmuOPZjxO0JhFvLtekPayDMPrX3STh3Z6HTb8UJQK8NIYfKQ2
bb/Km7twMTSEfkRuwgCtCiwCO+9uclzPKeRXt3b/5ibjB6ui6irCnv/P13lTqTB5
/3R4vV2HIv3fLv27nqFQZtdVDovPDZIfqvlA9RLJfmKbBlWiqCz50xh9i7pJA1f6
T2zwDcBS75ZAwta5utiUUhUTMFixnbDGRIrMzud1wngabCmqrpdn0jQR8sEbczYi
lEjJelM0nc3kKXeiOL8rA2WXvcxmG06j54wza7VnyZKxmx3uWJnTP0l3FTozitV+
OjFu4nRL2uh4ezQyHWOBaq2yl4lMGPRcjjKCiuv9GKo16l3zqcq2MvGvNeEKxed9
a+P0IbgH9CLt2VK5zzw8fZWHcsKAQcjzRS4RX3xBiuEtvwxT05oKwhkjaZrNnwhU
pZjYVnvj4mJNTBlJilM0IIUOkquaVHwnHKJG9ucAqY39SoWLCo7fqLgLtlzmsyDL
1LsGUxLPpXaZoRP+3t1AtwlThDwSXaz5kJrTXuzqe8ZsT+IbjqVA7MxEPEM/GZIc
tzYodrUwSZXB8fYgF1Whv3kOiI/2PW/auXqRYKZXsKRdFgV0ZB3HsBMDnC28uQg+
5lelu1haPTxcS5nug2aHiBWmFSYHDXrm/9LaWW6BgnkkkDsi5MCQBqdPJX3VCnU8
gUqK1nGK2TH9zVMb/o9+WXGe+elP2QzB6gsm89UqgtfnY3DdAzz9qcH5Vvby8fVL
n/szGitqh/8Sdr4j9oTdboZFIhg6LF9Oh1cNbGXk2cURMpoYd6h9oY/zN/q8xfeg
Kwp6b1FolzaIcucX2Yg/7Lxg5j1tQFg+qpROYk3yt61gUmg1lWXptNQCzILO+kNB
rE5QndjhDqWFW7+Ct8A84auKLQyoBmJ1ojxnZdAmeYNA28ujyu0jWFX/ezxDt/1e
0wHDZ2tenL8SRnx+hWDwftkPahci4JccFltvpC6Zv3yK5kxk8obXw4/xWHdHZUnX
fIaAGTYbrd529eXbBgtZ3h8MG/87FM+iFdZtvGPEovqZOiZNRdM//c0tqUDfAWmt
j5g6wpimXJgS3osqpcYfNcxzndSRRLs67mynoEpMlPTdXr3TdtJXVvQ3FvKCdFWK
INrZBZZ5J+IVMNMPFLw9DrNarXhzV5vkiZvLXEeIo4WUznewHiTlKfs8pRq8XMNL
eaE4EZgagTdjH54g4O1cHvdOTXBvK6OERJeymD2O8Ai4226cVvP/CAhaas7CMdR7
egMlpwifDmHnl8gBaTrEM3rYPC6nxravwWyVOJuD8LGsz7fBTqHJV392q3oKKpoR
filJs5iC9zMCeTPgVAMJMylOrxg5rnt0mHSYFx0UPKu0nN1WxaXN5KaqYUXkqnlm
c3+I+5dsvBWJ4JZHXHEd+FT0L9N7gOmeOlJ7VDo704Nbwkvka19uFWAt3BWEN8WE
J2wfFv2qVgYh1Ak3tjTLY0qnsjiCoNQjpGCc1/rmOVuwy1tsrIVmmOIJyYdKK0av
ZMM9euBcoxSjz7ik83xtjcOJgLbR6Zy0NEZp48pYj7T06LkR0pHQsWoHEVyLXDZB
bTwZen1wSu69cJpIVb86CtVtCXqTTb3sJ3//IkuQwwY5ouPPJuIZvtIkqfHYYnRo
9SBwQ4DPo4gekQZAO6PfDFq0dWJ8NWeq27p5FXl8O8A0+E1ttSv8EutBET7q7+si
9cdWYAEKNwqei4wTNebSYGMS/e8d2ZNE4sYxpUknl/0w1dMGVEpcuatLOz/U+CQ3
pfUBQ7+DPlZ1NBtU/zi1fNNnvShMV6Jpgs/38zY57n81+h2K4iIIdxy/LTiKIhed
oulM2D5FjhOc4Km6aPIlA4u8U9rJJFOucq2kPxdpLSCLHY8I0AnHRuaArrhJqyKs
QIZ+fc6Ry51091W3rIG8fXCGTMSxTNfFcJ8yvEAKgLeffu81Fr485/6/GmTg3N6U
btV16H6GzRjenUAuNHeYyFbtGpNksKiI7vMhMFQhtNgk/xJgRX4Ax4JdHXy9BnQw
K4cvHQFadBOqts3ywgHr16FlLPUYYXh92VYyYiLahtLogrsvVB1clwhsmGgxyBb4
gNCSrWBFPlnHlmzt68Ew0ZVr6XOESNBd4odnKRY5PLrRH+6N7jcYrWMLxdBwXy8T
mjuZVm/3UOmtkZ3thi0htOqDOe+nT3kJzpuJA/gM353+8eI1TtfNvlLgoL+8X8ju
XlzMb+lofah/DK2d71DgamFbIe1jEiffJkSRpkDpVz6dI6zm9lbHB6sSEIqiLuAr
7AQCXjS6giFpuHBmYbBUfj9Qhp1qIab7f54hVZvjEPle1wUDLaNjWgqJPwbWycZ/
Uiw+f+LBxaegnK8OBUmf3DKjsdUs20eZBuLjaxHk/EqYuVf4YHeEBmD3bCEDRECb
ruu6j8ug9Xh3dMnm7e0rGyUCpowHEuIk31N24rYX8PMHHfU9ydRMAQJZoRT8cEAJ
qXoMwuiIm38FHfuu0NJujPehSAZ0iFjC0KfXh6Y8zqzpLllxT2Bcv2NK/nmoKg59
FewSKrrcZOe3usLPnWlDmrC27cfBritAwGT6HDEzeKUi2dZro3ho8xzQQ0xJYRKR
Q7QoB2PCPPkDhTENTYlI8of5q+3b7Tf2BuFgfTFgvdYq9ZHPS8xB9G7CsVN97Hx3
g4PLGqBS57L4cy+zNgDqq+pgaLYqZhTlgM/xDzOgQjJQ4SI+pamC2eGZUiWow6mf
JNROA6q0Cntz2KthLvfIvv8Ov/XKnZE1WIrmUbB2tWYE80i9+j3kVFvgWsppRcjQ
WPFFTFS4ZJBesLfpZgTGIwhF2tdt8QL2mBqoVwOYErdMq+WA4m5/Ng/0b4GEXAJw
iRC/FzXj7vqI4hG0NUyc81/S8My6MmXa8mo36Vvo5OPMgmz7kTr9/btWvcIYcA/x
YhZnv1ht+tGfBOY2wJZ0A3uLGzwfpXs4JWLIhKhPzc/FF0iPLMrtFmoOVIfHl33V
pbd24vwx/drb02wXjinC7HfXc3rZwcYNTNtGVb/eTCggehFF+uwp74aQgBctX7J2
gvKF7d406FLpjEBlJJQu7ZeSgkVAHSSc928pVjlK6dO73W0rs9kxMYyIuA6KEm3z
ETrYDtvdFdXihH/ncviA0wtuKUJrM4ucQJFbqaLdSXZsQnZCJk19dmDtHbOkqDvs
8XjUOgpJEidAO7YcyOBXRGtVBCTxb53VIyknAqk7DXcaVTfs6Bh+BDeep72hDd4e
d5vma0GrV2s6ovQ/3VEymTvJGi1vm7243Vzsb/4aQDw06q17yQShdfmvxXIgV3An
WricDKyPSumwfbfuvQy4SlftYpf67AvUNjuR7dl8xXHMZMRCSGAC79cE5OWjjPnX
nWwycwxHcC8hvERI8BNlKQW1IjWkB2xQd58MAgRbgue9AxkDDOJ8Os7cymJfd0oA
lO0Ol1lbvyTU7PP2tPo/yzTaCE1JrZ5+MEAZNKax0dIOkTi42bFZCaKHmxaCMJ74
kMyMt9GgyDR4UZlOVqWJO4ag/PlJD11juRRr8hzHHzV+znj2p/Fs6ET3NUBrNHQp
iaPIamB0pAq3U3G+lXP/Pb1dBZa9IjlcjqXILtlX6RBvouxCDhdZLsQAULib6tA8
xoaqbsdxlrW8U36If+dW0mVnO9n8V67MgTzsjEPN4JtHrews0CJmIefRtAWg8ibv
KWpjNB/NFmIZJaGG1UOt3XVJDKxGAvAbayIhU7MSHrPM9K+I395TUEEkgIq/+pFb
CDDxR4UQRr2WqDAkPjLYE8ZRwfgM7Am+99z7WeEvxkSYZqFIH38BVV/LdqWBjuXg
F9k5SzUzCznCrJQeKp3c/DLNNNETkWOXjKnvzJh1QC6gBm5khtfZgt+AvefgD+zi
6Wb2X2p78Go97/XqIfw1LbgNz1uqD6DjA8xoZxeRv9uMUG1wzNjV0HDO9SpSIrz1
HaHuGLE5GSF0A/czcUd5YjXHsvVz3RhU/BRNSvAwyu2mTsMDG9v8Guh9jAT7bGgF
0lkhjZtY8IC8xWVvzHbj1XeioTCK/ANSyDFqbBUJR94+RiLzrdqWuyVUuDJmNdJu
IdX3vpOgUwOHTCEQG4/OgAk3Ub8xDXFWZAnGHordZeNvw7NMUAC8iev1HUp3hKY0
JScOwuGAZzQC2QYJyZ0+L0SwLGHs2HbgcUO+Imuc84LkkxnZu+s8cfMS4GSjaJPg
bLd0oResYw3n34igNofA+ONqTJU0g9LR/DLeJoQ0gptKLzk6v+xNil3hbZKmrg15
j7juAhy2wthwqHuMoe1yh7iTwdjelT6kHUqLQWdHz2OO+mb3tWIoWFCoxFIMw9vm
mvdNewNLlD4INOHzdkp5lF78e55OR1JjMpyk1r1Ed3Uhdz02N9iY0o5/K4YD6tE/
sEDMTG3vqobfV6NU3xaum+KrY1rmK0uhn7f3upzXci1/9XbmqyYFEUQrycKylgip
7zxYHCw2IWvZEur4SzR1U1wowKT9upTVbEcDnMwUrey0zzmUS7f8CqM2GhYSX2ER
pjUGecsPIQAt7X4tNXKwH7063ILF6Vspku4tt9Vrzfq7fsa2CzVrMgcIQn9LdYMn
ae5ObVK8Jz0EMv/MklhBB6c9HJFFkIJuSXweHTBO148Hib6ZiB06QGoVs3+Hjk+r
tOKzWqFwvNAkB4alOxuzrG+Hd7pu1zg8FDeKEiPeelOla2qUu2eRbOCQIL/PI0FF
e6TuG3cByFZFGbQhZg2UNTkO99YXiC+ggZ0xC0HToeug41Cj1qXcYVJZfISpHKzd
7R9quYMuZ8m82PHf/9IbtpI9oRwUwQ4Hm6JX4OjNSqlUUJW9L/miX/QUR/iNzJax
ulZzQ8jbpirDsZuAQTmM1uNTYJK/VkcWlBAVunajQhQXdMszsqH5gx/kPuMa3/6y
8GUxi3PVz5suKkW6p/aIxQLDcl5InhFEQ+x/rYCUuTy/LJqNOmwtFBVtlk5+qLnw
9vFuZb+ZX7SacF7CWfRyD7Elop/yY4Db7VpN+gz2Jntee+N66Xp14WSjxHb4OlAV
dc314kH40CSJvBuBarC/X2MthyNMamun8oh3FRUI/HbeKw9U/ZtfivSAESP4mIWD
8ioazPu5lNXLIFN8z7ZgGNZstlzphd2THnAjFNJOWELAI3hvqv0RwJ9G/AWPpJ2l
aNBJae+r3fMNODL8uRAGp6FmfstCPIVlg+bQ2mXzvCLsYxALgOYticAjCYhZMDt+
nfuG0zrr0lSaNliY6kh9iGZWvrI71Tn1LXQX0H2NxuELQR0bR9mtdVZu+Sj7JQve
TQy5T7EXjwfkRnk8F+/kG9GmTOnJdLQdIYvdgFDfg+Y7GqHbYEWRi0gGNvKYtESj
GuTg7KJpRY7Vx6t8uNdIob0fUErpUJMFj+n3cXwKReqsMKv40BUBBmWxHfzOVeC5
Y9nJmRSX3wzqB4VijfxFwepcQngO1okICq6w/aN9aI+sC2hesaMmHAe4/ooJ5qY3
FF+kcSDaHLihn+jbdR2RUbb2+kIMiQGhHMlF3Q6SkCX2DBM9cd3leNkfLhlVlQLe
XG1bUaRMHE/z/avZauG5IaPzMm/+hAXB/boAR0Xa5WF822MDxZxoHLkOTTJ61QLM
73ibtTOTcw5CYoPCMwknqz+mu4FCRB+ZW0DS7b8U0ZnI5BUx+J5HefJSITQeAWBV
tX68g4bOnEUQl2Wz1AMvxeuyURSW3cEQz8pA8jvO4KQKKdSSg/DMpG2gKoxLtFSn
Yqbs85rRhDh4HRcrE9QUForR2ELrE/RnwfpwcCGzWSYjdNtj6UUUhGZKmyCWHvpW
BQdAGRiKpJy+TKukUvDWwNa1IbSwoMTiBDtvFFubOUEoz9fPB40U0Sny2/RgyaR2
uBLp9D2kU4RSd32Ji8FllwtqU5DXo+p59nIxT6E99y8lprIZt/lzDIz/AqJggIyK
Ld0S0hO/E051qO+/Jrg/UL49iCwgL2MNakwzv26NVvqAN+qelIIdzbXD2ubAQ3qB
s4Sl0D2Ny7qQFE5z6B/RpsouFmgMbfGJy1Iv4c0bjQyJxohrlK6dr+7D3HThev8r
sts/C1re5OjEEn9kQ6fxiTN3DiqHegXkUBaPcj36h8pzs9njixYvXwjQw4eByYwi
aETTx49EnIlxPfS4J1rvvCpX4L4c+WEwCgg0mR313XNeyjlYNR79X6xQsVMTFzhF
4Vijk8WXhcJ/MLizYwcfI/LTheIVixa0bmXFs051Zdby5LHUmuj+QiuaeDdQxIlM
KSPICX/9FMAWDqHqWIHWJFLrKF4UZl5pNtf57nTbfEToMkTgESQ/MEyzwBaYgKX0
nHpbcvAqegnr/blfl0DlXiC8xqGF94AiwrQ7e8JHywn1jZkeIThkLzGIHZWGWu2V
QBeAD3EHQKA65u1vQC/jlHsCz04ndl2C/70MRIdE9XOFCVbK+VxJyp6XUtnj5pVB
Tx9X5pKMCVSjO1sdOYYtSJKrfF86FuFc3TLVXanDB/f5cQgKDHC8ZFjhLKZbHN4n
8HjD06IQEbB+cV7J0/8KqYKQRx5ubvXD94dXhHwlY/SjCDy+sNb/O59avmxk9SEg
TXrCs/Kmbi3qyYC+nb1haBo0MCM9AingowFcbakJtFk85ONrjzYHEb+D2N92Fxay
TZWx1iaaQyhyQOzBJ6NTNSJtLkn+KdFnreRrO9C4u8aMjLtln6JJmw673vIQZy5B
A8b2pLN2MNsdVW0BVuPBUhDc4nVt/WKFlYMgB/knyronvJpDNJxEDfygvxakXIuM
DdMCZyO85eKbBQC2mXdhdUklFncIUV+tpdWeRBGXHz6E/Zznxj03mB+D16N1ZvzL
qFn62J/F+kUyRWhDDq7dSWGNbRafV/ejh6E2TPa6Y/lzx1n7wkjDjp6h2G6ujVcn
zoZTQkzP+AXS2vueFcF5AqvUeF/kcl0vveGvh0rOa2RteTE4IH56aGB+ctCnO5wF
pZ3dH0gAtbcoXGt+0W7MANwj5BMs5FykwN2BIyXduD8lTNl0p9pPR6faMCoGuAOu
0o0O2NxQDc5yfOr4UVnZ3cl8ILpFv6OgTC3ZSe++74t6rel87X8Hk0UGlxAsu6lQ
LpHfi8yise+njba85ihoiggmRdTdwhJZdaBV3V9erC6ixqfIPRC3NPHB9xtWLhfY
IFZ2M/ZkttfnjYNey5VoSC/tazqxzS8IiGfoZsAOdDZXhjbC7eYBdgr8T1BCmNaE
46WcTtKoD9fsFHUrtkGaCmJVwDWHBjDyt2y6aezjFvU5UrZFdrz4XsSW5ULwjiPq
QbHEbzWrIJcckk5KoLYEmi/7EqDu1o7uiFEl7T+VaZKHv9RyT4spe18wi5eZ3OoS
kWSd/mvaO9Js6FIot7KU9it81cRMdJaNjyJzkSynZK7CnUWjH8cOrSoSk0slPxnf
we02ARr/KdDdBR9bqGZrXjWD9zte8k3F+PHI034+IXFdaCm077IrSr9LzlmgvgTs
xMdSP7epbGx9PzMQTYVKxJvKeXgHVmigWniIwiH+WEKqQAjByros8bysPKiNUli9
SnLvz7f7QCdVxq6zpePC63PThgloYmiK3v4h/9j1RrUjyatMd/UnnK4NauvY7jCa
OEV/SnOX40r/8+gH99qbxs6rfGpASvvt3jWWaoriS3KLCM0FkIuG35Y5Qo4Udmls
XH1wBgYN0eXVhGGcGfX8Vrc0EvVN5fTdHjIlKwEgqUFp6loaIqTn/ADeu6Z6+0FJ
itqagSVGnWrUuVek3cVgZ69Gum7gESnGccOGqj9yRXOseTH2UizE3hcLlby1CqJL
ojqS1no+GTAlHbbYghtFvuoJtfiafcYRQ9b2Y/BtMTqFu7GSRY9RwbF9Fl2THR3H
TZXlJXJVgZvZRvX5HmXHLUdjdAjkPY07BeI6ZaqRThzH6NPTXILx4PEEgQQmWcQw
nzgGyCaSQkifq5oQa3bnqmRRBWiaeUY506hO2yLCd4CGd2Ul7QQbLXOD6kHP+XiR
rrNnaDZhuhPW0q+h64D3zEKGfblRsHrhr+Qfj/RKo5A/Dp9YDhoXBTqNVWQgADcl
2wv1JTLMXZKk6dWL8Y7Dg8t6T1x5pc505MxlKpmKU3XfhA2mO3zfld3k1cefTiHC
XLpC2hLvtMOi0q9CINmr0cmffsV+xBfxR+CBwh9rWYbhfbaAUHBzb/qIiTiK35+D
dsqbxlomdl4IXl2IRpXglYs0z84jMa9J7ccceUUY0ac+FcR92aLSqCKgAlBcb3Nx
4z9CdYGz2wra4WddsuYnhhgnqtzNQgt+d3LUv1ghiNiUNve5+gp7jpo+7Sh6FHxk
BZ0vxeTyJzIaoOFZA1RKJOe+FEQM19T6+K1ZsLjqD+9yVwcDPg5DkEp9F1jB+ttc
1lL1HB65Q3mdV/XYM6acpEhRejhp80zMWvbNW7/fx9z/JRTi2kUwCFJ7smpz3Iuy
OCJodOkEI3wHtrMyzxpkgToaM2e5QdhVPlA5Slb1GhQTcDeIYr9OEcP6YL9bZJmb
sSqg4aIJnqeDvM0sfUSsI3sTCqFHqoAhvBwLHC2x2ipV8MvFyHMDdyE5V6GS/lQ2
bjhy2NxyYu1MfeUV/fJGu3qW3i1zVFaKoCLH27Ju5Apyk49f7fRtIYALFGbCCA5H
zUEV6FesQkGVyt5qoHbMzxuuc8boMzsdgrCsxNUZjRHXt++3zA0DmacI0O0jubY/
ImZJgtF+2kOY+bY1t0mcnE91+bZ5UnhgKgRylHLew7CNkKhFyZwI6nnGNkok/yUq
rz8b69rgxhASDXRcFKdpLxRs9M9WwYceEdAS2KiKsyCiRC3VCLN5M7OK/My0MypB
RpfNIXdsviPfLaSt00UzbtkVr9ypb+n6xlZ15mCmb62lv1nc4h2QODLjPb0O95RP
I2dOxwD22EBFbYR8X/cB7g2SdoLMBws1mv0HVkAzc3AlV0C/m2q6zHrjigOgHgg2
U6wfLFnSb8mkWQiSYjozvrgZ/hVxM+D3l4FGX3uXxpt9lw8yxOK6w8NIL3lA9BMp
lxwVsvM1bKPaMpmX7QBa2LOSeVrKG041FkbjZVWOXxiSOIIV9YMG68inLNznO474
P4MzUR+K2E62eC1RFpg2eRMCmiLUuA79Y0d4Ce5BkxzFlxg0FAkdrWnDSh3kqEbA
fDioxEJBiPh95GAbohbuGWzjA8c6dledsmFYqUUUtkYDhxnswgMYmS51gx2VGMx9
5+7V/iYPOfkpQKobipslZ/F1z5LXEf465ZMwPjXo5ggTDYMrZttBLJNgdbvgNn8e
Pr0rY+1kk9dyZdynloO/8Vg/dB5HNwrIpLNe+icbI7A9oi7Y7VonQPeLCzp+hAaU
J3ytAOgpuCB6ZgAMkyNW9LGcI7T4PVlfG5+tJyuhe1K1xYdrtNSAlB2GD8bxB5+E
6dBBEjEN9ScoP8n2RCGIi9d1kS0Xzh+yuu9+ozPi7Gq0px+xsOlx+JUm62paTVRX
E7hH2Z678FLcWbKIroOSvXfzfgjQLcJ5mcEIy8IzikWuCWrARflC49+D3/Yon4q8
QwMwh4zPd/dd4vGVQ1zyc3zBTxhWERHXl83Fa3Oli8b6VVZHFWzDK0azqx4grswR
Jc3oZXvaADJCEB0ljemTAQSf9H3z93KVdtX410Cajgdo82bQe+wu0w4HByMCcU3n
lha4IguKwuY+UAMaO/N1v4UaiHzMula4Vlv2u9Nsd6qAGucR7zcfmB/S1WG+mB+E
BUrj9ZmUq2yci9scoKlEwk1XcHkUyk9VspZkh2e1Np2tMior/vjKQENPNy6SjMA2
if4E5f+744kijzdYYi1Nalc6A+00zJ2hzMMcCznnDKE4KmRILQlpN2MhLW5EuOo6
gK3WQJxxFThxoA9f72VR4m1HedHxl6WGVJRm5VwnFJkXOk97f+NcimwXS95ALtTb
KNqhcxi8mBg9gok6qHLIpt30f3xE8mt2qpFQSKBXViszALdE50Qis0zvJhxVOjCh
6wQoKQykPtjf7znpRU6lr3lFOM7h63OwYLbpWr8DmOf741a9GnsztEz7X3CuBXF5
j+JTzYGqXr/mMtbs9FvebPmotOTOvYz6LVRJHoLA40xgmef2vQ45ZopcTN4ougyo
0SczD4SXtWxBYOQpXnNIqapT47phR+BrIrk0Frjhrn7JfmFigM4swFXEEo1BciyS
lCuYSeQZ7Fa49e7RWmAifjQCIY5iTLsMtO47ujSswyRFBGLYkymJCgXSyvVamGNC
LTNwRTx6Ns6B57/urfnlxHjaxNWgka5nx81GbI8rNxkBjwzf/fSdaVb86Gfaxkg+
DuY5Uu2czM1/x5IlXUgHX2IWw/RuxsRdUWtnCerH8srZHUek45XTj0B82h2K7Y7U
anpWxxClTVNWaEgSe5+iVL5GKOUznmnuDpUdpaUaAiSQdptr3PFtuUoqHPhJnfl0
qKwOHcFOIyqOlmT933xisKYu7cuyxNYcFOf9x9pioC8h3JEXxKtK2pqTJSrEyqxQ
nm34psuelbVnEVZPGpsq4ERgHUJb7hla8S0nQF3InHZ8VelZk0zOYzOXBR/dXc4y
JN7LzJ0Fl4kWq/iNJhAq1jRwRU6JTnIh74IVZ0BUAX/3cdwLpSk4Gf/cCk2U/G1O
iCvfUqsqsJX/vaycASlHp8yFZtDGxtX9tWzmEx2v1ltmJZfbNBOMLBy9SAVWnSAZ
nOX3mA07v3YKL0xD+GNAtl0cmntQrV2biIL7MDGMiypnzAWErktAiNqYcgY8wjip
psZXJhRFf5LIN1/tezWj0fhn7L9ef8ox6Nlr0xMTlD3yjYeJn0ONx6vbx5X+9FB4
rhQWHpoH7fD3sHtqmhfLcryQCamHs/ClHELsE3jmvApjBLHxNZPFxmsZgT5tsyw3
r0yTOQlL5KVQ2uKIT1MhPXVyUhJVSrGl1WW/7wOXKyy2VAEokBQamLspo2yG3n9n
B5IOdMAwmb1wN1wRrRc/xqUcbUwQK4heN7ejP3yon1CTbZ4HTSOulZl5KK5/pNWU
47PQV79RL9QftsOb5RlK2JFoxh7SWAMAWXTJn4tiqGxbVKhs3JXqyITrpcqwsoe1
sl12i0a2zZlwSBvrDBmS0twZzVFm548DlegTjxDSicnvAUxsXHGLYb24LN15LQ6S
jKVoEvgFmE0CRHH9wABc9WhOVeNEPwhQAh9MPRY2Fsz/5RryM+UeN0Q1I6Pz+Qto
n8r1ffUCzWo12WMvMtjR9S5Bx3ZIcQeeahVvGYXjimgbxfHbDsyNJbEgPXiAqnnd
1cUvigviSfQOZ6s51MTQxRuVpdJZF0rByYJAa337QFLfK10+j8VMLQRJafz1kg8S
oSqERMOfXvyOdC3s05gUcfV7mf2ntAoLPEvWEgzR7c1G26zHb0dsqGVzrIscVQdu
bXHVtslxIDyolakk0lSDO6T907NVHRQ6ZBw9c6jK1K5acI8KXHGS7A/8DLMWH9u0
LX76NCfFgfskWQfbmC44sAg3eXc7Sg56OdH+sz8qCB0kA0VFsQfCFCQLjzu8qlG5
uMjj3aPRQNrBsr9Y7L57zX2JrcbM40Gans3g4Z/zFN7e6X0Jhlc9Y+7oVXksw/ea
1ktktk3bqUwlZY9b3Hz2IAoJgrA0ZDZ39g/W7zjotTJB+MvefvmkXzxXh3Zhdgar
2yNGGq1+SxNa4LVhLhF2nRgu1tifXa703btv3/GK64P3LcOEk3a8ypW0CIWrryJk
k1+smQ6j/YjPUPWSwP29yawbsezsLTlAU7l2qXF7duGVIAHbYNDUfiPeIIlC6vjv
tUtylR5PPiyKyTWQvEXeDOq0JdulWFi7H3V7c9p0zTeMUVSo2/9F9GAv3iBjLeIF
GM03WrmvB+CG2Y5FlsdZLMZXbSj7xL2GpZ8MFpXbfJBN8khnYgHE3mc09KNNuCoP
egIaVPtGXTnzpKK4eX9blljKE6M1WAxlkav7EiJoUQC4fFmHigkSMslv7Du6Sk30
/hYNXa8TBgGlMS3TW3RwvCypn5/sGmO2k58nLqANwAmZIfMb1LpKKP5tdtMetO7O
h9dWQJy/ltwSYeOEqJj3Ewgc28XBhfIExRkWQVXxsXZ3T3NYQvwRIS5LDH0VzgFc
wqcqQ0Rw38jL7PsXP5iAg9x/60yeABczJ6w/SryzI0Ja6YFUNybfuVgISVAhB2CL
kw3k0LcsIVJmThIGlDD8dmP31IHnmIimkvVYtjkPNm1B1zGUvNeeaWpYneuc6t2R
nrRuqQmYloS/8DE1CSEUv2XGY1HiYyBLH4YrxvkANrIJJ5fmLMtLzEPbUwut8FvH
S1mPu6KDJTpc7RaAZj9hvAL/tHyjkN9Jtb7RcYs73n1HYGefdJkuDNfQEsd8Aqjm
f5jRLGknP1l9EJYBHl7bOxhDlHN1uWU7ZXbwg9yQk29c046nBcAt/NySKdZMP90S
pFoQ0wCReW4SOY/clfOqTGyRjSrbvY2ABpVfXkyHALmwQUyFx0ClRCsZxIPWkwtO
PUz5s5tdIBPML02LZAfPcFMn8rRtqpc6CK9bMiheAxE7Yh6lodr2eoBI7eKhLeQp
dpz456/zZC3hIiYTj3EAoNMLfAeHdpqo2nDo9fm8PqXsVRWtbuYRZox2PpIH8d1d
bhBKrg01otG2Yqgc+qcI7179imZpvZyeb7B7NRAdzkWQpx1USzqMovn3hCyqtcEE
jAyT7KYYvSKfTdZ0h0qPS3FvJMwKEp5+2zB8tS+JIsw3JkaTzKgl4s52tFmn87CR
iXboO7vIo0iSE7b/+F4dzNV61TKeywFlRWbbufHZyl8+Ss9gi4gPn0GfkrpTK6Ml
F45ciD3jUrWGo7ElJjSb9sqv3E8N9pn8QHgLtZ9p3K9eyOzpAtXRqP/ksCy/Ibkh
zZCvqeM9JkL/QfUM8LIe05wD4FDC9wpAPjRPWeD8jgo17RJYf/332SIjHcVgBB6j
lzrxL9/R3eMlGK+BH5Rocf/j7bPVx7mAB8uKJI4ooPpB7UNT01h6p1vEL9KJ0mf9
0YJGqGuB4CSemSVsh6m3psyImMfozCEQsyIPTMeQzNNvkOpDyrwI3TZFX4mim20n
lVwztAm0fYOVNf9/pzN48wAVEpKzS087H96SGbWPai4VsQ0Q4fK7WqQYqJYFFRsu
uqG6PpxkucdnTwxRvb9o2tgiwqo9QATiFAVQ3eXAkz7vZS0pMhfzLbKcltMTlzHc
j+4xWlIwCWOfReCYfSR1zYwANUC9TFpOIhcaRRt1muOPCMI/rqnf9VCFfl6/osVG
A8+yrcVeH63lBfHHXO6mZhsuQ1as7/GO+Q0e1Kzl4mKeY2oab+G77gjZdg/EcevR
cVqCTCdGuYrlrCZMSg5jJciTUE3VAt7i5KLTy6vfnaItLsh/+BbjH5Z7GmPzbpfp
RAGeKEQKj/CNYPRE7fuwjLu+s/JJBWudy4iMKgoumCUQg7gzKUwMznDmHcaqTq+x
0yH74mK/JTxJjRkBKz/wlr1DfdrIU3Yhm3/PJwVa47RtrlqlziKan1RyIVDzlQqN
bvKgf7L69wGmk3ARjVKh7wkszVn8O1gyEuTJVV9XoM0ISnfYUrHBVpZL9wv+PRpR
uADmN1bYttguIEKBoELuiOLyC6BGl4q9Kwdb75cGInccvGc17KuOj5dj9nVKXJ0q
PFklYZVai2E6FytohrHKTRLyM1WvVLl3hBeuYY4behvQ9N6W5asDlPtKmVEtgwHc
tKratKoquo2T8uGQwuzlCT4lnLL0cLY8F5A8e1xvzvrjmksFYIAQkfTwXAiTWKTA
I8Q5FCvIrU/5FBDS3Apnrkba2B8cwLqXB7fOUFqQJpYr1nohEIk79noSTnQAW4kt
R3HuYZm1wmBwhhPNdH57w1RHypxoXVoxv1CEj+mtFeXnHRBNm7DrGoEwlA7heJEg
9GeGx1RPg/I/rlzS/cMG2wFGv5NG3mqkZNFSe/0hpbhCqV/1A9pVF1oVoJiJxqeu
rPqO9pQKhmFThQCs6jQgRZv5GAAdTZlkT+slx9RZLWWjE2W92b85gPpID+lqbyWj
J+YP7jS1HBOZ5//pcOuiH4bE6lvBHhXoAsfjqIg6D+9tE7f3AOMnVD4ZzWN2vnD3
HmOeVXKkUFVcLooWCcF6Wq8NMl+DUueawXaSWNUhPMOM3ZA8vHxwrcRvPWdFZ0gN
Qc4Dnl2gKHz/nN9ZVOt9Axp2KKF9U6rrL+VakMJw16m0fWfqezOX0Ajmc7Es+/9u
B1AC2VvaQLpe3255EIrtKGVjIbvD/cStcCgZXQ3Ny/BxQtB/zsTLE+R7I9ECWtkJ
eL4PYsEbskXVfNYlDN8e97ObisXSGBH7fqiKo+C/YXkMn6/4Yn6zjF8/tp9Mbec9
YyALp00eo1c+SiBWfzuJfW7MKffP+ERP7m8+r5OLOgVH0kUVN42+4dlTPZMzgjyZ
12TMUPWcTAZamJVzsRGggfP5XM/2c7aqRGrrpKoddwehgG3nfK8GfZRdwapS4cfk
FncVqrKkcdFSJM5DcnIn5e6sQ1ja+4jyRE/I02DGalCnWIJXlSS8Ex68KjEgCaud
YjWOBJyfDZ/7+M4UgcBbGbhGzvQ204gAeW3/MUwGPNaTkWj7sDF5mBJlFio4Abmw
xdfoRPpwUMzCNWuwWsngCCsJjtV1P+T8usLuTUuK+CpSESviZFD3UaD85RYnjYpe
jBxXWD+L9ZR1S1SdGmgZntGWJukwTEjT3Rpl59aXnwo7nSOqPokPA46gIiOMG/QE
CyT4HJmF6icngP+JOhouF1XOdtPiq6j9E4IucVoMvYsLq6PfA720Ws3v/LwtuJzN
+3lK8DG8AE95UQHT7DIbTXArRfKWz4Qu0mOKxvze4/cbYfY33/IIW6RjlsGAeA2w
Egcc1cPVSodBKuCNAYfy0BXdafBRLr+mhM34RfyWfSmFAohf5j4FFtRj/1kCZE3W
4Ku7ifVafoG0jxjzgI8uGuMjrmF6aRfMiao0Cyn0DNwSAs+Pqe0RLtbJKaLIzC30
tbnJTKsxMsagOQvkKU63Dc18cBjcOKB+ra/VmauJw+ZsSBwtPDaXER7MgJwWAY2l
LqQ68ifPXwI4fQh/Nx3E1xTq5B4jkRxM7KdrD9HZviuWHKTAAXmTXqrjeUi2KlhE
+sHj6gkXMaEizW6ZNTO2C5zATT/+AKIBcGe4+mZ/pCxUoPaG4GP6MkwCoMraQz1I
9me3vQ3iN8FgHNRQUwNoU0TWZzKix4Q0j08giU3hVfzNP7bK+pMmKvJp5LpNk9w5
XEp86dXdBiG6kpq2Txm4SCAPfw00Nz+DbK27UzP4SPN/6f349+8573yaM0d4CgZg
aUcp8LoBHZ1cCYD1zwQIwa6pik86qVKO8co6oPsDHDf8gTeiH+gHnQe57NerMy0U
QKaR+1cE2sT/KEBu2t3Adl7Hzk2xYA3FaT0rL8f2ufF3578dSTUHLIe2yJC1aSmB
SWntL7SYSUF36jjNFKeFnAIeQ4HcOxIDuZhOttN7/qdNAyHYveX+QDco+UqixBSS
7e9cvYjjJIvsK+3CTas0ERIjrzwgRZr7omxjJKTBc8DxHl3Ue1V8pBcVaGKm0zIK
7vOBoRo+1f7+maFuLh80NJ0oos3yLo8X5ru82oex+IPE3EqZR+pPCQLnQtY0Bs0g
WHTErPcZf5+SZXlYdLqCm1+CHZP01oTlijVpOZxavfkJblJIeXU1VNgwKwoLIhmN
xPt9ZGf51TdxalX22OF8Wlj+1S+y9+qiRzT+TW3o09N0zoQbPfUCrDQkC+/W7/s5
a4NNjaXVu72obd3t6vsNx3sxgMwaPHKcezS7/5muVTd40ANxHm+9eJb+ENVV7Qam
p7iGXm3Bn8WsyHW85/S1MKX2aNo6bg8PLOoF1S0nyHWTDIhhB8WFZ6dFj6LJLBvL
/tPmXdJntLn2ItvXvY8jW9IfF7wc4YjyT5ZBM4IvUveMZ/6WB5JokMvFPNFpdsc1
Vumi/kF1/XPMWmKk7qW2PHcizv6Ki1AdYw8Zexy9kCxIkhw8fffd6M7Ug/Bk7ko7
GC7h5FRJ0PF+/hn1zL9qthAloNA9Z+xJDEbRCyu08rBDrMbHBEWWyBnDXyI8Y1ju
hfhTUnGeJ1CTwoLs2UcjbOG8/cOQqU0WXlcmdW2NmDdv31RebcjP4wyNsRswHKbS
ULcz8jPhV39N1SpGKE16K9NnCfrkHPhBMq2hco+KUP0/uNFRrLy/s1qzkx2Egosz
yYLd2iJ5bh2POGEUcLSCn00kATRCP4YNT7FwSunBF4SrbeuL+KmYAIllNqXNN/WI
EL0eX2apT75vLp5LFSLnu1qthbX3ApBvFE0HGzNR6MetuXotXHrMoF86BYc8up5V
e0YVd4v3PVTqwC8Km7IO92YS2oiib4cc1r+T5MaZSxO/JQC+qCyUTGHmokaNsunU
veIrVHu7LLwH6CC5eqoDYDcVqn2zm6DA4aFT3XS4L7GAIFCa2DUrwgYfG96uOHjM
rRH0ET9Cva5eHJ7+5apYpwGhwC4kwrUFXaB3AZPxFWAPHL6RZp3D3YysQdcBwpPO
mmhsak1Di4xOF3ENJkhpXxmGd4UJ9QQYUpR8AohigGnCWf2T4Nagic7RcxWx+6+O
/eKhvrmywnpzzQ/Jxy3ekeAulw8n6o8v40QTnZjmTkR7MkIRiaMpJH7SkP3u82k9
Z22h672lnsuL6jScbsjqObu3LmsVJ5buKXDhEX4Aiam81YhpZvlg+up1rw+WGxsJ
8wnSyCjLI8FqOTB2mZ5/DC1KMwr+Ob62CavFI/at+8ha+YzaRiOTwrO18QeniJkQ
j+Iu5xzBc4wLyR6Vlh2clK4pgao2pbonsbSvLbCsEUOnNR0Prtexcn3VLLzGrOnG
LNnRYbi50KC2IGSUoze0ulK2410Yn8+x2dNFXxC2/YEZy69itVeKF8mUqz3W6ejD
emV+7j99uzm9TMfcc/75ldX9NOSkLv33HDfCZpKskX2Ec17rHmBNQfa1dDg64sU7
QuEj9pfqRqRHpYrtCBEnqiCbJMn0ERNHWvfuZZnSDfA8+amwkxmNVEonD1fB5ehb
lckDEAy41YcCMT9AIkAlL/iT+yhj/poKdd4X93brj4ulM7lxDw4u4wxtyoIIvqc0
Nt+t8KHesgqhnH+wndGzV9STpngxf3fj2o9tPnTamFLMOlG2N53PuakmkhFKfA4t
mzHwFSZzprZ4JmIYKRRw0mN5lMKI5zFc338qJTqzE+J2qgzd4+ATtFmzz8Mqm+QI
D7s6CTJ7YWGaB8K2suPqZMmVtuzPF+YdFnta+ayzV8XKcLHOzVwfVtKBDFo2838L
gNwkYNi+08uirLM2BpbKrMmLNXzJvr+uu+WzTxm56Hx7J7oMdAb0fRIl20whXF/m
5iArssrB96RPtyBtsV2dzKKO5X6Juxk5RI1W2+HWdybk69UiHS5rRJm4c63TSg29
BYtXFz0exP+Zszono93W6Uc43s8Gpri70T6P4836VBAU7UJYTiubdCQnJi8fHSp+
ZHZlbQj8fpwAefbLMC+MYAw0kCIa1Kzo+GoZrJSLqkbTHNOKNo0+TFEw8PyZkZBR
5XE/rkm+ZRORctmN1Dcs4y3QNIpdFmyYPXFdtdtpx+ol3imYw0B9ci+T5hGaYX5f
r4RU8sfZiCbv/yjaVXI8g1T37zSOYnbBY6WU7ket1XFDjiokQ62wA6F9HSCfkcoE
KDJKR/NE8a2+8jm4qKWNKQy4UcocC9dDuF4A0rg6rqvPkcKtb4j5RRuvRS/HBtTb
/YrNqLAW9eV5nQw1LYwAUXmN8B6O8thot7QEM3FepQj1M94gsuNVkTlreFDo40FV
mf8OG7wuYm0BpcWOCm8yWs9AsXZQT8z/66RIrhGml1BSjQcucrijzPEHLYvAiu1e
LihjClwDByoBudbaHeGPK7FPwu4c9fID1n7+VYG4G3/EhxQSmN2ZCaLiC4ULjlnO
vukAh0CsYUgnmvtDwXDIL/d7E46vVIwHhtM013oO+dJmngycYFw31FuQX9jxuKC4
xrTOso/q2bv8s6yYnKskylNeZUtnC5R86bRMSfcffmUYozuDkqApQmVmMdF4ZyPk
bYS7H5CEfU19D1Fzyxp5AECDoe2Xw7zETH3hskC+oiOSN82xpr5ASrFe3IMrFjl/
WVlQ5h0WE+rLaesXTY0tnwaA1w/zkMc0esb5EqqJAt0F/nBgauvCczqEN6tdedSt
d6/UZ0gw/W+SERGOIgXc6CGT5MWQW1Gi9JKHgyQeK1tMSywDRF1Nl6bQCY14sJCa
CO4n7WFO02L14RmO3TCJ3MfNRzTvU3//EEhZiAEmRjzjxh6oEXu2iRrhAjPrGm5B
bZ27RGuNF7cCbcUBZrlusvOoS2pSPbIn0R8LBbxT7HmD/zmxKCeVgJ4riqS19Cs1
bgEbMEoN/rhCPt+NF++JMG1xMe9GTWjBU3og7fJ00NAmJgKWOT23llT2b18mdQy+
At3u5GtOtbXmuYncmHIL6NXXvmZ6q3yA5IkW1GKdDIdsa0hJgdgbonAMs1wcDtBk
2CyIJe0IubRoPiQOBJg4ZZSukH2ECPvXSXYaRfuw8D5BZLy4pLTxfc13UiH4fgEJ
3+58Bu/iyfm5SmoFKueAr2xgfo74q4NjG1pJL95SFuAotX0bq1y4vJXpElfxwc1J
Pf1ZAT0bZB/Chzg7GxdJVOem0bFTLOPKGTJAwdCAziOB9My/8xGoQmpRWx9K00a6
ZpxQd0gxiMVgnynVRXJqYmzdAjRoIZbQWe0W9b2mn8FVOJWdDXs9INT3WdwexCgj
gqVoV7LwpNuimpO9s8XCX3TTDnzS8A8XahdO3TX0VzSV178ghB8OJsECnyGZ8NN2
rlvBg2SsZX4R1RiI/UoJchc/tW4BC93cu0egyj2xJRm36ALd8+vaBbSE6J5Pb7Pg
ZVTsbJsl/BeTUdWdXwc7AhTPGbD+zIOaqWp6wFjwdphKAt/oGfiEKTPcDYD/HiE8
ocPr634lYc4gwSHP7wPsW/7u80YLUO3AFO/Fj4QawdZQUC1LeCiIy1ER2ysvnpGG
fBW/8rMZ9IYfRYeAjRb+pmvLO03fwMtIdAiS+1g3uoY+6ierRinCM5jS+axXWkX4
clGTJ0aANnXyF0jXsSSLp28dQ1DdSKxI9UGvE/4Ug93KsEItlclSVWDsvnWF8KmJ
Gm6K3WW4wm4dQ8RskG2IxwS1/U6b6xAu5/8ZeWRj/XXUhTpdZfpG7beT6yaDsn1l
LmGS5ZC4AMzo74NxOW36r3wwpO/l3BV4ZBzfiz8ct/WvP3b1Lo+oKvF65QVUsDMT
5JBPOu2mjIXZQMw61r50J9FJ/VedryenGrG8QyK0SGM1mCbStsYm1eylfIrC3WpZ
pPFHsKziXpiQI1kRMw83fe4YhtGUAmttl2QgK4IfguCgS6dG47TTfkudD7jBJNsa
Sk/AAFWwHK+vkGD2h2oIFwjwgsYMbsOty9EpAGOHVRRhj0iCY52kPPn/3LFrwXly
7iN+z60oMp7QXtFfkYAiZpgzkgSzMLsOkkwUVGJFvndMy4mR5eKVu0j2ZNwV8xZ3
nY0UUa7yZab6qBAF4PylgRyckoSZUZf9R4tscks6ksnpz81PEWHvlm2NFznR+mJv
YgUh8wWCyITFObvpDUECDJl6Wz0kDLdYDcm/hTB8jo/FSjLJgdDoW2rjgPa0E4Hq
byB8HID5gxMYHOw/Uc8so+rVnRn/VkBWd+EpOwFFWUvov7VLx+GcgzjskdvWaTQA
tm/Y3t4F+VMVr7RKYmpPTeR6e5umnkNyhiUpdRYRFxoU06aRM/lzZhvy1Sn2X6+q
VBWnbUDv50qHEgci2vWDCWJxlI/844j7qrcGkMG+YkV9ZbD4bBZz775is+5H+dZS
Sq7AzGxHq+RLwlLSfvOTw2DZfYCE3J3IjZiIik24RiuR+m2X1ZejADuXXMtyYozc
o6sONZ4HkBfHojmhbq9MskRK/my25Kb5tWX2GmhqhKfD4xTNIlfjzUhrbqSmbVS6
3+S4m/5bJ3I98TRw6XAIesxz7F5wGywvYpa9X5ToQZNGAtszdvC4liRcNu9lokF8
T+fFwR5fyRtpodkkN+hJnebCTsJuV1+wcv9qyp/MwxmJD0TorxKdZqDya8tladBx
hBzWkP3zP3e2UGrVo8kTwO3RMgzjTAJr6IWexwtLJby/VAxoZG7g6cuJJ1iwl7HF
yDGhGqtgB8pXb51pWFNuKimljOHsgFa7ZiiEc8AXnoK2EsNk3vEnxOPbOaERhUAv
I82H/7PyBpl1rIBAGUMa13pixepXdPeB1epoKG1wP6hJncEp6C1IqoFQHEmEUeOa
YCIToKHkMWw3eYxynSZI6uMDMh0IzEuCmc29PctM24vbHsMRgEIkZAUUYR8bIYJp
mjoKcdk2mSyb92aYQgvERPKMRoLvaVnPOgXxvOUjcEAXGkr9atjoHFHJm3N9suXG
SaH1AyJROjWiE4vd0kSexC2ZqpJpKSO1C4OPnVa9RtbXFnGx8hypEZhY+iRHCr2X
jCqcVmzqLvUaHWQEoeFlQhpZxf4y/LdTdsCbyS57b676ahzccHuFOlWJ3AlnhjKY
HXtI07hZyiNeAjiFJik48L8s9l63kyBRnSmsRb6iV5bw6xtNsSTjVN/DBAhiLrrV
VkXISX5dfyDHw5yssethmcpdAAnUKDay6yZtRHu3j6c1hUQI7K139gOGCt8oGHwg
3TrrIJ8mE1HNy2g+g1RlIzcTebN4TAPZym67YVzUrnjsNvFa6vJzyxnfJUW+EaqV
aHdBQGJiE2HJoD0S+NV5bOSRlfEePUaZJRrzY6shYmDov9DLq4Rj7HljNlcBYwM4
mHLckMs5u/zBPiU1gxcFU6LC5vv2xN5wtSKoZMecPrZt2tyAdE4PKvTpYbFGUvBT
dqhEiYqe8Pk7VyuO/V9iUAKIlP9GAa79gsTmtJ3Fc5MEXIYW7eeg8NGzPLUY0uvw
FCP7wESa/bgMOoH5wVLejbHyla5L9TnlJYJLsk6oD8pT27S8j4XxgfmcVXYLnYLZ
LoQmLK0zXj9fU3wXvBNhRcqIx4OablUvLkhMMKFP1JSK+ojlu7pfKIaE0WqMHI/s
MBJPEtzcBG7uz83WzfZke22lr/6zvPaXQ3pCtKSHmD4vos2R4yDd67N4pg44Kz7X
JTOqyGiY3gUHiMuGq+4peG+VvQLm91MkEJ+qyv65hAagQ2JyX5S4U5XiGyOrbS38
I1irExaNIJcWvYOeJHfnjPNTEtH2kkUHXgoJqYaKA98azcbRtz76u77sqqY6pLQ+
ybgVQScMdbvWOTeMGYnp9f2SlqZ5eb/dOTsjbqbJ1ria6V1IsSoapyXydgfpQtU6
+t7BJm2Z5cjcE7T/N0eCOAE0lRBt9DdLZLNDkfozM0Z/JpeidDJXCEBK/wgWh4zV
w1RBn1r4X/WEcyg4Lg9MhJ6RfBZ0aXVX2X/XuySgupPdd8916XzlprzI2E5Hvzmg
MQvE4kDnmDEBD3xDFYZyGyXzq1rlMkQSZfYoYBXyjEgunKz/nYWhFbkSARSllwu4
ftnqjhuikLXgwpFuRgX4TD1da2yXV0hQjpotKwXK/aPx4EoPEfCbTwl5tteqHIoc
uNmgmTifWPwF51uJnJzglR07/6DQ5DBH/+m6GMpWKAgXDMP+NW6MFpMBkItOCehE
dLXU6HOxnV6B9wT89PVQBNYYvCo/WtsLPMX74Iy64g2FW+9jFFsZgIxEO05CRCDs
OB4W9dNWdzjlMcJhnUAbijKygTW0uHn4JhRIaNkam/mSNHucZFdy25/OSUyw+uGv
L5tB1hfa/TykF1ODZ3qpL5zhB5TUhM4VzeKl/9IMsJ2mzxV3sPa0qUh3nfw6jlW2
QUrVYLVfbskhHaN2kahLoJkRjf+4KRkHiaGOwO2lnqJd34pLJrNEu3QUmLeqaVK2
3UR/yQxEePAhYd4jvr/RVfQ6byOsbbo8pLJzObUSMRZtWl5OqU2GbsSIC2YMMz0E
r3VkoES5iNXgO/4W9bxRuuZ/HxZsUlL0qp6iSpZFpspzbrkUIJcrfrhg8+erxgLy
lJGXjFiGR+EWwDnj1bCMG9w5ginzu+l5othNrfpFYPnwdPJU/m6cK2D3ozLcakrm
NiRv995ERhmZ2bWY+0/zwHX5iaAgiuCr29gYnywu3TI7/hHMlkyECO5BNgIDaWT8
lXzRG8uM+ZWal500YhHEnO3MvtsUz45aNmKH3PM8uMRW3XZj/4L572BBWY5I8s3m
QsNmHUSpY9HDRjUdYxrHRO4/En/Wh/F/8GKXrSkMAA5uolzsUINCpnwU7mt7BJW4
CFH30AqWZQtmG3/w83UBONp0ODUwrmzZHTJHODJpDtF7SjOqrDht7vENmrcNCACa
7tzyILnekPfzGv2oTwcRo9m1uSydNsk0Xq5XCdPtREX/u6vdDLMHwhEg1tRdFEbZ
5yLiWq+fL0kOWlcq8c2iRjit0YvB4iFKwaNx85hBTkhW6wRPx2XnRkgBWM80kjNl
Q7s5WNHrKCbjkslvht6anSTpzBM8Pp07DGynB6sIxSc5c9yggSIjYHPjhOr+ehyL
4ejYj1f15TXjyOguDELYd6V8SIUwFSvfOe9Pa/nHCdubFVfX0fZFBo8Roq1Augq5
SzLLwhFFGnbYRHUDPZ7Ue/uDVS4n/a/hkJFxeincJsPaU0au73vMXyIjtCy10eSA
1MGo+E4RnMeHrH+oK0LUyIT3mWrpEXdg2wHLNrywmR8F+QYhp8OoWHBqgcQidb5a
PlRhZaY2uMS+sqk20uMYAgf9PCZRkHidrMmTACZqvZ/CEF3HDmpqzh9JU+iXMyPT
cSzP0jcBiBay0Si6KEcfK1R7QUiKudEXUuIe4q23mJ+tmhO2gRLhoZ5yWxjdlnjA
MCwYJQp646HtDXBqBoxeS+asS3e7PRcbbGbz7CYfqneCUq6s0UiUn+SKg3HKVg0s
wuvyS5bIM3T7JtYnwk2ZBY5e5XoAQZq4GkGJ1Gm9ZLesCnIHXteZwnQObGnT+4Ow
p8FFf6jsY1m0F+R2MGIRhP4ExsDe67kimHebbiZIve4FtLqh1zylavho0LSFpzVj
xU+KOX7gpCSHrDxQlZf7QWNa1CKOwFvINBcNA0IavkFz4WU4m4RAirH4Yy6HAaMB
2X4Y6zjpyaHkeFp+qEELlkS4GEuyRjvqvaZW9uCL7AzNPGcI4hrY3AHAKuBmQeyv
vpvuQmQ6BTVsfR5we+oV5YI3x53NvXNzeQW5YwpnS9Lefuw/doUYEtBt9hbqUwMP
pqT6tWXHDYFm7A1OJi/DJdv4+86W2rOjSwskQy1lLS/JkkdpAoOOVf0zg4ymGf3A
K0d2X7OUm6Ivto+8ohlngrQlH5uId6nCfwjSBfbJHNm64IHOvpaKh9l8TNwNT6eZ
1YyONhZphNao94hyaE7/rF9P6+XmC4yNxkgeiQqZYQ77xJA3W5OHh/ChefcoO1TJ
7KIyS+rhi4FevSY79xPCMJ8EK+AbQUZUwsuyBQ37joI+p1xCEGesqyXL4e1OB+vy
Tjo8M7sg5M/o7dQL669K7plWOzAioC/7E5PRgHSstRqS5th7bpVJ8Y8gV8Yft4Md
9vpeZY1b6W+nCuf0IAZra2Dh8mVUAdl+kpUE3VVpZPhjE53Zskg0F9lqlk4FifkM
xrE2mY4Hj21SKYyyZ4FhDKArYS7ZEm0Hz7bsPd0/w/pvEljhI9hsA0Cl1ZtYDrm9
ZBC9dGPfStlsGbf0nDrLMcxH9/c48Rq/oELA/Uc5BClzwTXrBf06C5cawmXZGDbl
SJTbo0RDuExXUP9JnzHVxUiwv21njtx3cEUnYeUVOeyTeAQSvNwDPlYCnoCK3sMM
nbPmxHxWhI2WcIeJ++oLMj1ZSZAKPUDtVkKlx+rsBoJU4r2oe6lRJxvScqarcRBp
dr6cWMubsLK0r9+NCX8ZwhFyZLXtoIFtjtuWOJCTfOx6KHfJHE9Zd0bPZimhnM/3
XD/uNhWWXn277LUftJbzGlrnzyYsKD4zS4uBzAFw9uKPm3oG0pLnlHin//PiYiKx
afCNa8aHQgiWohVG0wSNSqtRr/nw4xJb61UucP5HragEpR7F3ueyATHCG0EPexjw
gF0k1hE0Ypd5PgDW+Waupl2EwTB5qel+uo6CU5vN6zlMG3VAoLivoW2ID5bYONj7
wo9Tb9iAVGchaX0vbS/LIGHX6Jr4bjoBZlmlVLBfEnDDVL5esFzBnuwC/BWV/tH8
e/WvaG8YmwzIEPFP7ZQSSFD9/QLXTlIqM6pnITeAeBKmu1TchZeHPBGwoVp1xfyp
OeksoEgl20jkpymyADooN7BtojGAXw6wOJ8s7L16495UZXY8PaC2fu0VJWKHD700
NEuQxSNqRaQsra7ZXW2l6qnxz+xdSo4BHIXQp1mNbSBOP2n6XAToXWpvd72vS474
Q/5PXEFulJMH5hjgTIkmunr2pz/I6pPxP4k4+EVErlq58gDm9sc+0aqX7hj8k8z6
EgC8C5ZgAGdAugf6QRN6XLnePM9ne/T1LyYzwCJSmRPf9GDn/fr54h0pXJaOPLMi
3ILOmdmgtMQGh/ChiaGbOu1nZK3dqkAYvkcajMfcWREiyDDHFhTygd32V7X3orX+
zhFNJCyDtyraI13n+s2kK/8a/WULIHmlZfE9ixvOPsUBEeyj4TujyWyPiWtZosDk
F7q1SP5FjCL/amdDMYuxrVORcfNMcOYjEMWQmmcqsA/KtSD/+m3uFtUUqRFe8QUR
nlVz07frABpuAkrfVcpFP/Wtvb4TUSOc8kfLJV85tMkKUDt4BFg0SZp3C1i4yf/Q
nv4JVr5SUMoQ3seqbiqHT2zp+4iP/UJsKBYMY5V7+76TnnJIPKlhKwdeMml04qQt
zvWUueJ/Fnk8O75eAYOh3Oql8ec1kXtyKX1S4WD3OwfAn5IfEWlGP9X3WA5AWpPQ
6L8pSKV3RssFKaWEv9Acx77CL7WxszZWUGVxnxQBtU3NR9DuxWFB+RkPYoUCJlh7
S9PDNJdR+eWVeYuHBzjbxSU+lTBT5k+CXoRnk3z2RTZRuhMkA8g6tm/f1l+FFR0X
SCu7bhdVWJOjevMpXDqVJ5GJlFgvgS9YE7uIJjwKSr3lSSUozP57lyfIkR9+D6GX
cea/JFsjB2snVP7hsHQYjCxj6/+P5TLywjAVwPtQ25AVmshiGhAt30FVB9vCbZuN
3OGyqMgU28G5GyqDdG73IT1ai3mteUBgTkiyXRuIBr3j7wdljPNV2559XbCowssx
wZN2U11EW9AGT0kYVJIkDGCLpWNYVRrmj+ooHqlX9aUr4pa/LBlW1AtYTqu5ErSA
NZm8fejevWgofGbg3ZiCt+wZPt8BJKvQt5XP4WxGqyGxYU2ei32DXUJsTLC+G1ee
DAPzji3zlnzUgFNWPe80SGzo5ZwWz6wXBx7zY54gKnzxEIU3/PkqAxx1nnBYOmrg
9SERwziOm3Qcb9agbfdEOatpq7VJ7oqsp4wTCYpntjiaDZ0oebFv64UKaIKmXJHU
I7A7Nj4aBEW4QdcNl0toNfg8FPwmLPbDiS9VWDIFoPwgu9/vK9MkSyzpUw9F6uLQ
4yX/4BkWKODNRESj1PTy+l+8QAkmBqdwz/nEVNAGeRzhxAmD2Qn62AA3kszRtJQ1
UNL5v3ddvd6wnw8C6ca/DYfz1BU/EvTOP53fFojvlujzK1OktBRvnLcBKVInbxmg
8CiQOQIUxqXAnCtvESJCJQPX+tQnA+VmI6P/WVvPZHKjKiVm+E2FE74xWm0lSo5I
v12qoAe03L4pAJB0htYUoqTyCqWj2JLHFwk43ZJWLiPocrhhsatIeHYe5XJqJxuG
LVO5Jocs3g/liB1C+ARGE9MWEhYYDqfsbJIwms+lrn75qJBNe1D70KTeM0ycJzZZ
ImdI1WC/aLrA8CwIlrIHAqgw4oszUz9h/0G3qhtpw0EbEGo7pg90/Z5gdEOmLRa/
jtb5aDS7sdcHTzqTDpm7Xj+RETnaZCUFG2hWTp5ibV2PhHzJV1dgNK2l3sLHY+VR
KOtA3nWOa+fb6A5KAV255sFqyiNoAA4y0LQ9JjWEpRhaKy+H5bLcLIOiwUFnbaWV
hsys2b4Qw7dTHRztxPRGeP6oCxAr8L5QWjrIhcx7l5JOd7ivnOkFcyITbOesZxXA
pdObl53QLrDXVq+4mv5a5GaIWZbI8/GAYvWOWD0EriGF4OfK+XCnbIYQLHQJ6drF
VlJbLrmTAwjcbqO66VjRj0R4q0Vk/lrJj85f3REXgCbKAVu1jLZUkENw6ekXhu9h
J1UTOjJWdEHITiSm54Ay838iv/k6coJpNMAyoY2ye5aYgM6DAkxc99Sf05QGBnwk
JHvc/UhMwVMRSzSdivE+tFodYh1IzsSd3BgA248jkpo2QxlRozIet0LnjWk5lN7J
Bp1jcuhv2lBu+/TnEIP3P1oS/OddHDXfyYOwAGieCk5zkOMOaqTl1314mb0VO8Sw
uTDSwtNwE13cGUKexw6qnSn2tmktpCu0OYySvR9guy4h6Qb5/ZYEHhnobizYIOqb
ssNTlu8kWBuRxHS38WS0Qis4YumnuBdgFIqdU7BcJYGzLDDCDjEt/dBRnlbd0yFT
H7GATX3S/90BM2rbYptK/PabNL1nTBPAhGr87iKFQUkcCzAMjxc8VNCSy6JOnvmr
XMijwoPDZWuOGShczAhrt/TqezKDo8y5sntkhAOdot/S1ucjsJ/23waT/qHjdhyT
4UhwqrtSokeW8yRzYiRba2vbM4Op8uWy3yovqfgR2KzUZP9waA2zsM/HMCS/5IB5
B3oXNBHK2B3z+da0hi1zyz0PPjrSCfJwuv9fKZV1Yxftqg74mrNXcl3aMNSIBMew
2r4AvfCdjYSfz1YNqCSt0PDaCB2FZrY3L7XG5mqVyelzSmruNP7TjOhCxISXt2HB
WTbWA3torhEpTA/EBvPDyQxV7YZvsWHY+qMdyrQaQKu6gkQKu8oQZPcBkEwvBw27
NxZexK0mKzAlCzN+PRitQgBiseJfxu1gEVNjOncH648+sA1fAlhsFgFpMW3ojBLG
gZ6JKPVsHR1i2pzSbJZacc0l8nZh+re+AVTyQxuF7DOrVg9bsu6xaVmIfw+YcmCC
n+92yAvpCfgE2KBjQolCKOHj1GX3kip1+6QNyLw2uJGghvkJMs7oSiCRk4JJLqoY
Jyy6F0X3Y9QCZE8ZB1Vv1ux+o27ylVwpcv72Ha+iGNRe4ZeIW29ynkam0LBBuHta
dVx+QV/HpOjPycfZDGU7fg2L38rKTSdPMzya1C40tTruJhIontJVJK1r5vj7uGX3
+UZNDcLNeVuc8+basKmYx/v7AEYO8nDjuwD/IKz/B1acRnn3yLt8QbUyE/6WlVKo
SyMBL+p+58FcyKSfQ7lkNJchU4pJ1yybZLax2zKoj+jEPryiM30d/01O2+kCUduz
tPqNfx9Wzhem3tGc+jXP3+wxnND/SNX348fgdQ0hfeJfPsg5wHGyFsARsLqKpYMa
1XNE/opkyvPJoIqGx+IQdx9RqS07QNFKDvSIlD81mGm/JSvDJPYsyLvHcoVpZtp8
dsy23HdwIC8EVHuJH9bZB7cTeqVk5ZrBycEtfqPTFbLlFMQhUV7tLOFRM9nFa1Zv
DsC8LXG/kAfJJ0ZQaYE3Bwqh+HC274wkwr62HfCZ6PFncCj5NELdutL84fypcc7A
SLt/XNAkJ3b44/8utIsShtgV+3SapS6GPPhX0kisRF+OFAX4I23Qwft/MZbRVWOc
jBHl+POgZdKzQt+DC1ayQ8WWdy9DMWAeNCgdawsc/sBpWU8LDehSm7cAFlI+ISeq
kOdWsAGt8fvIRymnZFLsPL6mGAEBJcAsaUKDpR4J8tLXE0NZgPxypoZ8XrTKNJqz
4Ag6riw94r6zFMY6MuOhqxlz0emE46DDgnJDLq1m9M2NOu+S8Oo5HFHl0tCihHUE
nVaCjYKmk7ac4t6agGbZrdRlBzDWeMMAtU6JXXKIkfvJdySRKGxX79+krV91K7/2
b38nc9FRIOtmFB3w/kgfHnYUFCYPWhf2AzwP7fIS+4ib/+JtjNFdxvkw2BLf7CVb
gy7KdRyW4FeVTMH8SNyvz3FbSFJiQxW90aSB0mDm56fFJV8iZEse7C55QbOhzn8P
HYOroX/sBebc5cH/Mkma+jY81lsMSoDmGAoC1SnLA/31lLOOkV2HIVmznx0h1G1G
XYODWG9BNJvbBQjxynvxbFFkgNsUDN2beTCZI/r/yuOGUDZBqI91WSeEC/bXtFKN
XsgTB1dvAgCxIdtYCXu4n+mlGsdlle9kiSAOie3lEDvd+fTaR/lLbvyegRbvg/DX
TmszMCuOi5e+Frl53keO4IZNmU+0cG/T3UljMsXwjPDhmWcUn3sXdgyiO/Yr/Mps
ngZBhcgtq0wggQ07zeN6wAhdEZTcGa9Sk8Xdge+n4Xq8wHoXARdwFIItondupq6B
8l9nUUzbyJGDiCTtQ2bs5B8ymKDy8T/0R0HSqABg1jE06hwza3gzPFOj99JGEz9z
A/U8HKQGaVpSUPjv/5hoMgVmqbQScmIK6+qtZQ0w2Uiv8KjqL0ELxBnPKMwaps8U
fIX/tPrUnqNvtdFO1ce6vaXK036DMC1OYDBzSL4u/sM3vOs8726oBW0FtrccfpaK
W6cNrw3uhkheQIdiJUlypxjH64weYkSXGhdPC89nIWDKsj6PPOZvFJ3KCKippDHr
xyN3hh2GIslLHk3o/YTrzWgtRWooLdk7J++FngwMR7vAT0lLx2lrp1ruBObrH9Q+
f8qScSs+EpYX1N9MfKrLxRtSovxMxb2p8jfvwUZGzdPrkcATF9+2KVLk6CaWim8l
A4HUN1/2y1kS35LmUCZO8S6vlaeGoQB89INFIkxhoFbKqtmfIJc0abhI91tFY84m
U88bitHuS+2qV4A898aG4R1vN8zlH9H0BDsTWZNRl86QKGDjyPCk55jZpNcfSZcC
GMZXQlS4Mr+r4q/mTYNwRMAm3TuBckzzzrN6HtYIRgb4evCqMgome13n7CXJAjc+
60GzVZ8cdWVA6e8D8R4fHPCOwr675/1tS3xUETW6rwtE1Em13DviTTLVyQm4dldJ
2lZVVYg6QNk7i3E18vz5MzJyfx4h1DOUxB2BfuWIbhRK5mPStAuEeBj8Rc1OEywa
OeyZh/Hvk4PARXr9el56gu+ODJzq+QBZdSQDxcrhjcrU9kzq1NifFYXJ5xH2VwI9
ptY8a3BmTRQfsflXvfllteYekyvrannbNdJsTq9p/mifOkFgJuEzGeN2jhXUetGC
wYYsqDnp75M2LYsfPoVdQgGnZLXdhimCEwK21+CMJMq4jNo96Rarw2ejRppFqldj
DKqFBBtqFq5oczDynDDKOLaqTEcnCYYilLccARXnqsRRc8AtExFUH8pIChALky/w
OWipbq0yDvbbytBXi5/tmGDUbBd0MwIlY600LpzWjM9rCQUhAFNJ0UwxsJ7FV6NB
SHpIZZjsUs6Dkwhlyw8dBBhCio7aTNUZn0MlJpuFuE6GPqaie53VB+hScoXj0+J4
edqjtm2hgqRUIDzCEurVac0SUbRBNMe7sJ7xM+D4pcB4YDLUI7e78SLAVzausy2F
dlVXFcMVoxhnWZkrbF7YQhOK2HKZ4Hfl53GW0w9fLHZLz/VdVFgdBgY0HwYsJ0GF
rW7rBY873AD7CUU12kQzywPiRaI78T2TfZhAR7uf6z1moHlnzUsy0ivgoHqQbgMp
T7zUqg3PQhceKWvR23zKf5/ZhKtcGdM3FyectYuNPXzeyRZvb2Mu1dzc7Y6OcNej
VJsnLy1UdWJLyEuic2MP9GQCRyrXkHJ4CHVqmHbIQbLl0u5t5w7N3/BTouHtQkDN
XKgrPDZ0BaWv5u+kRS14vRdLUF8vyrTTPwLMNHulT8D2oNAh5/bbdAqyOk4ScA05
h+BVOyHmdGOe41ozLlF4T0yl3d94clew7YkWBbIlnIasbyjOP6P6X4qzJsPIKDdL
5u9YotRS3ar6f+Su2tsMSZ6YwfJeSQlgdflukZsg5ztKlCI+yKokFn5XhA3/7hfU
UaQgR85x2YDqh9pLEYEJJ4TAH4AF7L631lpaQWUZ5REYcxd6JU9gcZgPE3DaeVSp
1wkWyLVsVJKQ6dKMb4oRHYI/6hYukSMe5P3PiDByoL1ZtWEJTGbn2pyARzcehbG4
M5/ojzc0u2klaphJaatz06MsbxOvmOb8eK9ziAWnuAGFDHpDNHnVE4bapi9wCoJU
bXnJR1jDjxN6d3x8qFCquVshVacunrGbwrFWgXfM72tWikDpkiwsYliAb8DMkoaX
+iuYFX8tyVZRMqaEgb7NKnycwJoOqtJiLxKsTGABZ7fjiBAe+9gcp4agsnNroqd5
/axKZYWcJtxN03EfLUfgcJgAZPAV2TRFWVDjthir+S9QXJec7E5XkfuIHTWHYGln
R1J1bUUqcleXS8u0zFsvsprAaLChX7lOJK+1eNAjKFbI9h8bGDOfeIKblO35/L2h
Nsbw9XQDzb6Xw1GGxswWMzkL4Rr29J+VebfbbbQSNd/IunqRYm8GgsVG5zjxArQ7
Lxv1ZJnH+lecHs0l7xynSs9xah1vGNQ7jEeFY3k0a1k7G8Ng58j6sntN39X80zB8
Qum5ESU+ItBhrjTcMpfC6l9DE3dKKOHjE1S6UHie3BoBRSD74pt9ku7g7mN7O6m3
isu3+TuXW71za86KA298TWy7atxletXVAJL73GAGSe9D6y2uqt07bWByFlpOUc26
FkHL2cAiylvEIk3bugxBC5PbITJWUxaB+avw0lrNOncq58F6198Etw3DKTAcaLei
421/o3LqeWlf7Bflrq75yUPrLGQA5ZLBCP/5VSxawObWZG1meEGjLtrwBSSvX4v1
gXwAr4qV6w8l6rXPrAz7RNjzGoqnvK9otqCMp1OA6ZYYmyoms5XkvMqP1O2lbCIh
CJ5zNvd3kkww0TFiC5DYvcGRwGOzwI2AxK4Y9axlIQ6XH+0JaJQ+JgcjDBHJuu2D
98mX28L5hWZ7lkbBqe8Aib9r/SlqWPjlbXAiTjcV7zk0AcbalTbe0BXGraBy58fN
ql134IALIXdVFJLko0TIC0Sgomcf0KjQIw/+lQAcSle0sR0BpYCqcSxEBK3Oedwk
pJE+BJ0s29pEK8wAD1Y3neXLDCKD4NvjJnS6CfFmerYzDt8DnO9ZXtJIE5PCB6FB
tmXba3dyT9gnL0l0gLM3pzzxA1UodfXOmbeJBsnu6FEsE2re6yI1KnVB36S0Dsps
U/HCHuCYgfHqODwpRZhK+XZP0C2/8xKtT+r/ICDMyfXlEjYxOOZdxVXu76BWvXNO
bbQxSLadSh1PXL178ZoFEKIV0aG7Y+TLi0WlKSeZGY2gw8ArlQ2pRAIYMwmaCTSq
TMhS12RCGHeQpIr0hev3JN9QPdHTc1Grnhnd94g1mcg4w980PyR8TmFC5P1kWuFO
jY4rPtfrJVE2CZcxv2PJS3U+jxLcZ26s9BSg+4aeglQdr8gOrfRoGsorgu97XSt/
flR5RxVnQ3vbO1K7YqYwsD6pRT1TCU6DqsfmJT+LhrXAwlJCP1OWBQc2CkS++7OO
5c4yh1p21ayPRjugzaWMXA3FtSSKbyYHhXmgEBsbbfSBUPhp+sIA4QqKqncPQNVK
K5ruu0E0StfU3G5QEaDXU7JsR6sOSnXLHl1dvoq4aluuXXhUlHBEL42FOMRDI1vj
EcuYK29BY0SxkyKZ8DzJdDVXwjDtZfBJXjp+T3azHK5aV4+QJVj+QY5Y0Ba970Qh
dEIwEMpd6iBZu+08WMTKVyjQhFq7FRT6nqZ1PJykCqgj8M4/8lqh793mCJtSIhd3
Q71pNGh8rXIijOD2/rEA8SCDkhwnqzEhfUnVCsy4z2GSd12D/le1n4mocJ6P7QeA
wDSknkHplBJw34Pjwr1RdL9UTvlxCRbrj6WPwYpr/7hpneIXAR3FDNcZBlCeAE8h
vHvf4pvYQaWUK1ExSPiLn84lFbkf8qZaDdJOMVlYTgARWSVfFzUZ0akAiOiTdgCS
TkWtlxE6D1IJvk+z+B3I0DvlT5XHZzrZPCJWZG1p4eaZum8Jpu5RrYC26mEhVDBS
wDlLjnd+HBrthFIYe/cxSHfWcSXuP5MjDNHc2RmTfEea19833WNkQ+DvZKzEf/ZB
YhnQfbol4IFEW74VJJLUcBL+LLTs3rLdlP5D0Dz1/AqQBhMGqv1DBfDGcp3epl8b
NZvsuY/SkYY7bn2Lx6sHcV5Jg1DBMSVPf2nl3rkOGsWwWbsMAw9v+3onIdbItiHP
vtnF2KuhTA7Rpb1Jwmn+/ehy2XMGeVANN2l0+9Khyk9vkxNdsryaASL0O0Fqv7vb
OlQRf9hVE7P2Bz2s32m7a4/Z+XHctkltknFNDZM09KZcpfrBCrlK/AdxV5DfQ5CQ
FBjMBjwHp69KOJvVkIEoe2QYxqmDHvek25z0BsgPp/CJXxRu5gGCwcNg+qc6zdWS
OLONEegRA+a+JlqivpO19qCQBtxLW1V/J5jWWuanOehJupHBicGRR+sZB2CiWLPS
q2a72Wp0WHRJFw0mrBCYxODHX9Z6CY9yr0SShPk8X3vUdKvw2Y0ofNOylb6H0OUU
lnTO+u2e7kf/RV86mCG02Tq0XzIKWEp+5oIE5UVlIfzdvoS4u3t+8WYlG3+A/C8l
d7QFirhw6u1Un65Fvr7NLYEhA+PKYCanQdgMUZjd3DeGRGQhmrW+GL7nrmnfhUOD
8snhT0MEai1QhFoxVmLyXPsz9zls0iXVrEnUvwrEIiqdJsZciCq5GH72Z/v6wYAr
Wm3uNRXG1wsao78QqP6iKFW8yLVhUwXxkKxSc3CNMPvRJxzVaQiE9OQTuNPdFKcN
TYwgUOL++6RJ8uYEX7KxIKqImReTf1Vr9UaLkSMmdzri0f6TjS3OGapAXlO6BPGu
JGKhnCbGYgmgqr00KcZE53lMUn6L/FcYnlDUsc09o4XIZcohtEQFbnxJw/eHWiI8
lQGXPqXMYh29Y6oHyxaX3gRW0cUSFM4Z+YN11TvR2H9dDvrnLZSfFVDqQqpn624p
hDwa/UYPTaFh/fk7QaJ5nkrFKQ8xDze1D4LCOd/2gAY1Hu11sioVfOFdbaL2zfUB
/LOWl/RTuqpM6DtT78D0RPRJzGXbc11ruxTDUTm31v0ml+M1FVbgFJqg8fS7aYpm
O1Rvjmf5Kfb8kJ9A7Zd4E04ngs9iofwy6rCUZEonDo2mj1Fzh3LFetOfZqZOfRdW
jHujJqGSAZXhP+GbJuNLBevnShpuFvNHFEDVZXjGDTJW/+CYl4djMOl0asZyhR3x
FeM6lJ4/iEV4BsOjPHq799wqksvq6h7QGeEJGQM5ofhZZPJk4D4Ord4ZREhm3b0f
pZiDIitwx59RkdrUp3sF6MDo+HHJFCv2FizJFhX7dJv322Wpc0HRb2ZDHpS5FmPg
uD38uzKcykZ+KWxY4kRYblmpT08SgHbm7EjzIe+FN44LT710j0lbXwBDvfxKjX27
RuCccBSF8gwo+kjeTfMt9WKshFm2GnAQd4yA+h0c1WPeIIfqbkQZp6CTHpXN4y9W
IFrx9TThrvq7BuG1LAg8a7K/+e2uO9Ny5ALSSOSXcup1qIM2dWXoLJtg6LLUBsHA
MxtMBRlUi4o2xtaQgglmoS1N3SDv2vG5iSkGqBcom3mhVASfYBH4OPzkVrPiEUrv
yoqw9FqUWaTcJ0wGdMzvL6CTGDQM/rzWVIhBSMikJiH9mrBbga0AlfHmfNcSpPBF
jgkYGES8BOS1pMcnapdsrWsoHtKz/v6Myz37ykRUv1ob+SN1wjij9yflbTITJo2A
RMm2pjv/TA2BeGO0/Lk4U7K03EJcfzFDcAQMH5+7LlrwZdyRqqzNr+TZELEzeNR9
417MdTiS6YiqZAFoR/w49jMUS3+i1fJ7fCmDLP0fu8p1GYw9/hAF9wZoCWBUEaJ7
qDqjPUBai2b8Mgm0wBr3wSaryOuhRZBJRgU5+lpwK7oi8tX48rZ1Hn15ZIYJEK3P
YYYEG08jIO6XXc+osui0CMeFcmjoQQT8EsXO7nEy33ARyt07Mzhogz/IHiGyJ8vz
jaIOkIiJr3lzMZpxufr3D8qcefhmi+k0y2X0d7wqbO6SyhHc8PohU7K5nm6H9L1s
QDrkns4nEhwGNuGGmXujF+m8ZEVjFu2iNaS3Z/8+MOBfF0a8YmNM9R4Lm9Gtojwc
I0A++DpfCTMo0Ri8K+L+Jp2aq/s+msTaJlZfHsqG4O5A6NdU49gXN/VUBxjxZfKb
3YwdVFK+xAwThVGm6AF2cEy8oy49T/UCHtrwjl4g2H+4hngQA1Rhb0VZqv9U1rPa
gkV6TC1p+TkkNOP5z1AMpUcHC6gtr2oMsQURVlRKHI4CPtegpm+4A7/EqPUNgu1h
9YRg6DPYU3ngWPFuR4u9VSXriAY1zG4pwkrSl2jmQ0VtjVTr9XYBGHBf12xh4CiR
nKYsaGBkw2tRPHZiYk47slpuUOYgLF+XIuikO3nxgiYpBVeuitY9nbsKO/jR+doP
vTW1NTojhekHDFIOY4LpP5rgOra6owE7bmcoM2fS5nZKP4ByThvz2XbHOdYC5Kst
4sRFkdBRwzbEtRBysUr5DTd2NEdjjZN7gfKq/j0YLx24/U4qosUIRTVHpD7W7Bp+
f2O08d1lxO8iOUs0Krb+dheiRNsi7mmwLBN5jfBU8TprMjDmRK51CojrpbDSpO2g
jSJTqKkZHbETcZKaFpEhrf9mR5S4/WQtJhDF92UeUyxtJv0y070YecH0f854n59u
h6v/WTmiVXpj6vkcO1T+l1TjAXFiwVFgQNnMH42VmA4Xr1YSFrbxvrYsJWotyPmN
20TYxD93ynpllkJpmuPevEYbjY4G3SUGZYi7gQfh2+SeUrVvHXY4C1VSgW6s6uwH
Dq7rmuTtxQlzfYSYQTyigztj29tSopmTgTYRrQa602DncY9yfBaXoYH1uhqnizxl
+xospEKQhohu9qeiZnPa78E3CXJdWDaD5ivCqTGS7809YrxvbDm0RiUljdx/O/lN
tI4qOWdqZh9efJjiEmByeIAhruY4AmolsTe7k08zqFPyYBg7a25qs9QfPKZhxeha
tsoK4edic/EAbbionVpJIHFY6WheF7+RCgcAWNVlAcBz2Zh4Sm1iWtDPvWgE9+8N
tVizK2UAGQ+J7tEUGtLByt36JHcPUpjYHCrEYgQP926v3Hyn/FamAIT7UGpSczAv
DiBJiWowiVwWSAR45T/TJc6Xyd9xenfL3QX2/cdTYopKXbfvJti9GlX2WNWESrGi
5kp8HTLFoMFllNPBOeinTnbecxHpfUGHAefWEN9l+njj2ktCZwRjmxPumCUGmB9O
hRQf4VcaX7canRQ0rUVIO2PVluc/DZaEEYHc8i+VFaI769Na132d6ZnTW+FMWavr
kbgyhEwzUgC8l4OsiZYWdQ01anoLmyLa3CORvkZXpBjYg8bDqrA0jnVstvf5JZJv
RgchdT+xOuMN4nF3aPhTLL6vptOuBKqsyGvpC7IFKNxjL/Hm5JhTldrlF59PFOF6
TtHamCoyktDpnGh17GgYkc1VYvGpmRhcvKCH6r+j0Jc9opR9gWMP++7uU6JXXmgl
w6a5LMpRPk7QRTNfSp3zkbTXhxlZUSIhbx4K1QJckD7d737RPvxqhdty8Xku/5BK
AdvJKL7GHAf7niYnpXF0Gx3lNXMUwQB3aykLC6GW26gYpTF2dHyAVhH0upvgWD6y
HmfPvyjCcW0w2dIvjNo5OM6XJihqIp751ch5QrZjd6xMtNM2sN7K4sVpHdzO4THG
He7Vqre1QTAR9vBjrTSz/ZNLWioRFDu5OczB0k/znpxGS1sP1ULxU+iCmoP+yoQI
wvSZF7WROBcsFYdxDFYBKE70phzB/OY9kAtBQ91B+n8T9f9ryVsNzwT5WNv8I9wI
gTTYeHn7IPcJq144rPS/zQI3SRHyv5rL/q3I5fjzvHmT1EoNfC0q/C2Xr1YAbU+5
+JXOT4hhFm8x0ejFl2V0cv8RILBF6x0zbNMbBRChx1aDCz4hOg9oaDA51lOQYwFz
R26+0Pz0/XBbBVL7kaakcZi2n0+3Lglb7vdi7XQyI+F7IrASodoFQMfb9BnSZC0R
2Meb4GMLTTA3haUHY1o1fOA88ioUz1df52PCj+veX37/tO/kHZtep8mq2L+4DQmJ
RKcYi/QV1f8w6j78RyKte6S6LWZIu9FFCFPXupbTN+89hB8u5hmSvehyUHGyvIOs
kYGpBM3MBSucj/EIZG3fC5AGHjUDRDbN63eSYB+3cUmUNZOys6FLZZmC/andaobw
pOivr851BTuKEz/oYO5ie3khAE+kdSbGdzTM6DDpY7DgjBNdzycCzCeYhj9togjM
ZGdzQpCowQN1t2Qh6bd0AUDW7CivohGEQP+tYxtekcSDOFmj0+7JWp6TpsvUb0QD
TwtE9fSBN+Ub749L3LjGPxuEyxneQv1s+xsLXYxbXuzIXCl1b0xlJ21x6A9jgHfH
PRGVMF8tfMVNCsCsS26jT5vuLs5mF2bDOWFR/exHisCdCWuk2JD6BIfZjuz1rt9K
342n0cUZbsT1WdVl5i+bdvdSg3Rv/g4cm9dtNoKqweGwDjFvXRNmIWJYvYT1GFso
/iIMCoQRoPwguS5gMplO6Wbf+AUZdE6tXYnZRmBZ14X6+m0ATlYvzOFSmxD4g9Y5
G/liYcLkZ/mCiQfhHlrt0n3e178sv8/XaoAy79Wkfp/t2OiB6ZzCKsK/jV3cPU/U
d7o/MjgEUEd2NuKyG/M2LiFxmWFkQW1HEnulO727N2U+9KK94UOO0wIDXo5nRRyo
RAqGwRLM6dX5Ttj4H2SOKgGfWg3SBI5YncR6Q4JbBeMZdyzMIrJ7AI/dkbwMWGsa
rCq+wqj3LJzbbabfFz6pkpPZO30NkImpq/feHebc4G86pRzTCtqzVbY3IUaGJhOC
sCnDr2zfkaQcy9HDoRxuoRAOvvKwXO4f/c19iRhUxW7Eg+XPwsm1Ctv4X4RCpo6I
ixmjjSZ5AA0vxg4yAey5+5/TRcQwNuYhRUWOoqVWCVSFibpIM1yibf/QH372V7z0
/XLD99FUVoiaAqlReUIsoo9jV9PDmoBml2l8vJp//ZY3rQ2DHygsxjyfnsh10zBy
dP9vJTvlaT3C2n0wYCKxwy0z+yN7VF7vX6fVijyeL9asmAEnOfr0V0BYoyKGbBOu
wIxWzJVser6u0yBD+j3MAeu9MqpS/qskoryXYQjOhyCJzSl2FaaV5mIHChw6IW/y
XZ2ZCPrcsj3W+0diLDznnHvVK/erkC7urnPtxNBBsS35pHa4cwv+sPhwaKx34LTD
CuksbWJ7AF07QRw5ovAPYu1RsbgmY+gQKSdeH5/qKwzXFGJWtJEu0qNYok+uyQFZ
+EkrTzNyHimmILV62nZ5WB3SUdoUrvbTDqxQjdq1IgWtTJQ5Y7R3jtuu2YcAVoAx
nNoQjig92LVPndWdwGbdQZ9gUuDdgdhvf+t6kFefa1n+6P0ZZVJBQUz3U6/4KAkC
LFS46JqrVJuf90JgrsUh/Ab73knXLAow8id65Rhg/296Iye8dGu1W1Kc89wVa+ur
WgNakrIDWXr8dMBolnN3mFaxcJ9icsokRtK96Od3Gn4G/VhjVPSecxfCkd+qYqet
fLwXZvn5uSewP51gXDy2kBpF2EZsB4tbNRHG04VEFWvu5tcAKX9BGgjQBXaJyGV+
ww39VH+pdLoeg5tG3K+dORUG1TaVuYc3cwQnm+m7RlpAqrdTcss9FECjAda04FVN
EBbxSHbroFqNW2JxkfRSZJsH+oZSNAiDFIUoKKY4pE7oMSLkcKHWS9YTpQS2sAu/
VI70GOIpCXylUDE9LY4XlNdfB506FjkThBvMP7k+KxzRA984UyqcUQrrqmcVXcYW
V9x7yDFt3wYP5IN5ZA4DM9H9fXqHEjMZk4UKqkbMleGur261uU8vEer/vms/e/pI
ee2BFLpI2QawjtwKWduPk9SgsdANWDvJETehvE0Sz6SP1gWKJ+cc3KlnJ/FmJiRr
IkghIOGjr9Snl4SCASU2CLQtDJiebBUZOpZFi2zKVX0V5Tipg2d6dUAYSvT9fL4B
EXHOU0RQlIS7FPENTHAb+Bobj2GmhGJQM5eKhpoqvCEqrpfXSRQVQPNFJi2uolG8
wXEiZdscYZvvWV1NoYw0e6IWzcOcY9WJwxE2qphaxhmZDtLMLnsylf1n/ZlnuJEf
85qcRWC8cj6R98qJrGY7nUxmnv+Q1fce2rTw2mItrcNk6L1SpmQ+tTedqELgWkyv
JmaGHHGZPcgodq0MW6Mn1Bnbu0kc0eQ3zoxlHfGyjWENhjeUfJnuY0MtvS/zzrxk
C84RvotQEaCZsSoebP2z0ZAV/UcCR/kKnrMob1tuTPoSkMzSsG+dRGM/WQ6jKAvz
hMUD9+JEmth9WS58lOlNXNzY9Kfubnw/CnaWTXzdKcKYUSMcUjrS7uIISPNLOMP7
tAQIhUPkE1KBRLfjpLbZAneUISg755BmBmPX+oH8O7pSH158rKfwTxI6MSZvRype
XgkX/z29jzuvUAC7FzxuteOYbZanihqzcAoA7zQ191+kThwBj9gg6MwEW2fN39+/
EP2mIxyFH87AiLL4oJng3lhzCMGqH1jNjVwrOAkWO0umYwlkyuKNI5lwiviONg2i
0IBvAtOZphvlxsteT45CqyeAbOmJfnvR8gVrUITEyT/QGOBg1x7F3Lorg8whO4oT
CrT/h4HzUmj+Z+mxAsvne6zyCrt9BHuBvNIlRSlIKSI+scJzVF7KA3QzQ5Krtxyj
sasvdsS3uFMQHDbVHzD62um7aBm2dT0GRaSiVDJ3WqmYEIpjQ/EOWAsKZ272jh3K
MmFZNLiSJNijLairKMnu3e8uja8T4RSh2Y+HVXnp4GDtGagfKvHsyijAD/9V6Gur
e4GrWTA7M9VONfayYmUSfoseOA8iPaFYi/4IMueGiccNgTmBYgWvSYEIvPVNMqW7
XNiU1Yb/mYIGbvita/QI5md0oW2TTxxndC/ffYcL1wHm+k2ZNFHMwRFY351nbJrm
3gB0j2icvmAiVfWUTqdXldZRITtusUT8m8+27dLJ1cUQ6a05Quxn243q4NbkhvnQ
9PwjyxyCE0/0a8z5q3PghRLRTl7712O4QytGpPH3NdQck4rhfAsHM4R0aonw/gMF
6r+xu1CUi/2JMKDAAwe1VnigHyPmsRZnvY9fP9m64Njb8k0HsX9jZOtg26sHCFmy
rwU5lgViOXecHpStFzR3QiVSXgHrV80lrZ8XgIu/2XpUbKG94Bvw7mdHg7AyQIk/
kEHlysKVn6V1PzVJYhpUtItYEe5pzKGLZP99SYrCrDJJpcZd7GQAagpygPIcHqPo
Fwe1L3rRXFisy6TLAIe/M2CfQMKx8hmQ6E+FB5/klxkFJQbInuP2t8bha9x4JaYp
BeAKW/asYwfe85wtqQ+Nzkx1XU1Qo3iTBBltQMnMPluTfRf1Lr4WZyTvVsS71qDE
yLSEJD+lVSnZlJy5yJuzQIm+Z1Fl8j3pGJIB4NrxqPcS7Rddlu5i5pAzzufTel5+
jy6Jx0wkUy7fqbbKsmCrI7CVfts8TS15eMa1439sgZztQUGYggiV9q4Jyhw/+5wq
2HrjXZ1oVxDmTbK0aZuZuqNCXSg7OGEfvr930dwsjwZ0Q6vbZrMdCCGBLwn3uYBS
GvD6D++gdoJs/AEJZvwQeH22Z3CU/xOcANQGn49PixzG6gjQpK24qaLT2foBRH+V
QEXs9f1Y7R2gl9BM9ZNpWFF+PpR2jQMgDIjW1JQfp+/ublWO/U1Rs1QaCHSrm6a0
/pvS+v5mZ9JsrK25kclceCVshNllsgzY748C7VXWrSedpDl88XDTTF1Zd7IkSIOn
w3hpUHvbx9iDOIvI1vEpwOvWTKQy+CRCJdRp5jat8ZvD8LEERsdOY6p9TT1u8RT9
+rnAqQSGDLCM9xLFu58cBayNELWGB5j0Qka5dTK/PutOu2+iVt7SelABpTZG0d7H
UqsU+gtdZ9KQgPgyfDtzRFgeY2UNvhG7MeAHM4QJl8DXGVu7KFDH/JVYG/unJS7U
zA//2FY2Uysdoh2kMEs6fPcAbNHFaA3xzAw4TDX9GAvfN4+vaT+Pguo6nmzRjGXA
d8BGo4KavfKEjB0DP0U1sZ1hGujnLYSUBP6B5XM66mqYwFjU6uvX208/nnkJDyty
/KOH0XyPrx5J+5YBB66xxQckRTHUndxq6xVfxnV3VXKWOh+K9SdWesFVfXs8GCaK
fOsWqRp5QspvMD9gFSJ3b7kecWxvXo+4WsuYgDvx+AvmBJib0v798iWQRM6CVRp8
vjr2mQfKaoq869yRFu0wiOcnrKuI4fD9pIUC2dWrPjUsYy8FVxO8dsfvHRMUzLG7
5NLVqmBqQohurUK8+Ncrz6SXTyp95uNJhhMaOjvwEo6d2HlLcCIndHAxbBhkMvy1
YNWYpaXUYPxVUm5rX0PmKQRca167cGPgItjyZNWUwG+fNiycyx7CL08Ov8/Si/BN
KgCm8QLltHij54lXQHGFJR7R/o39QqJCw95dwRmAW6AoY1NKl+3lHs62fBiDNK2R
VYBv6/WJMKuvtO3UCHZ5qGRiGD+DlWNFyXDvsbogysomV43MGmJ64bM7o+xLmfvJ
0AZ1dwpvFkc8thlqEKcOgHOLVfNZUxDxvgR6HwJWhyV4NvKADQY3aWDZOH73F3Z6
yCKoZcP7PcEtn1nUbJws4FwZ/JD7MYSL0H/Wz8Q4LPWJMcGYnxmuoTAFfG7WMfdc
UAY9DardOUAdtCpvkRNYUXBB7l7GQwsCXZOI1KvPG6i5yEELWLAB+hZMPcccBlDD
0t/nX4Nu3tjvSXBK3bIQNmvnI2/0uVEpYGg/2HyNAyNj27YIGjXL2KP/4nEtiili
dF690e5kz+q/Ckov2jjX0GZerlpj/s0H9GhijZ9Zot5rwLp2Jx8Y0plsjOPSHjNl
W1xm8pfjyjhu9m81CiOO8kk5k8Z5mn44KPeIOi8DyBaJAPUHyHt2e1cCy9RHd60Z
G6ybdtdU0d5PPgWeZzNafXCuMREgixHolezNQG+R5lMd++eAge1gesULgy2tPsvU
9I5JC/wAxLuoUlk8sHR3g5pZFzHiyHvdmXvEQ7dgCWaIreTao87PHn9WR+7u/SDg
7joFdrUKG+qS53ggjROsaKuHE3TY0OlfvWFs6jOv9gWPdPc1NFUXuRYscWgiSnBA
BJhGIjeSVR+lsYLaMT9HcbxI7ukj+zreS71jRTfXQImTtKAMmPXa/AemOBSafZnI
eF9zxM2o6IKlzSZ7X+n1FI0kajsMGjg7xWIdUPJkBbVPog2Brhph8ackc1Ey8tl5
rLuCdrrMdYoRxuMP0NvsJR71SCwT2t8PZBsgdayMfYYYewzX9myF7yeSlbv8Mqu8
mARf4lYqNnJ4r2UAql+ueZaPjoVU7AF+ThtYmIteekoih/Xa/t/1DfVBZoynVIv/
pegICHYvRH0VPokaXJkjQILr0UrGY+HTd/IDf5rFTimLvsr52iLH4sphrRcmZIUc
ASIeAOd1SJ8zk7czUPIYOUALwWr/yu2iIEiHRVxW+qDsnp/yNQRFbCWR+e9awIfK
SE3JzTex414V8lOQ9rCwXyT7mHwfYGgdO0ZqWZrostMXufDEKxpt8HZpqTgDHkxD
lJTmQTuIyBbayKO3eJDHYuokJz6owObM0Bi75Zl6cPRngHQNgHmDk59rKvO1OrKv
S4yADjJQLxpaUbdoOwHxuaEUyJveAk8/SeU3U0gpUcJp2dn/5E7XySXC7sAbgiug
cQ7y47zmujxBapfjsb2F1TV08yhVnXFP61tVIoHQQvSAUs0aD7FSPScHdhcO5XU+
FUnkBDse2JDi2IwnVJ+6CEigYko1WuG2sIu9otoAHOjjXyW6s6/NhGzHVhZyLF0p
0VKEsAYj4VhW1EzTVDQL32BHsebiYrG8vcJEIQukxfM6+1vGp3BvKQCe2tBvMv9r
LFbJL3sgzAVJYSWM4ZEh65/+GG7WAf4GHaP27SLKyJt8g3U1YZtfN5Sq/v5BGQta
sFG326D4Y2spEZ1z6YGcxErBWlnFV2MilAs1uHUCJewH2j6XLWcCcGX3/6W4Rbri
lPCNvgyIBlAZXNAn8dI8H9dLfPZ7QbDoi2iWBBx7lTFXDjFeuPccBSPy+IHSaplO
cYUH2Qy5WTUxr1vgkaYKarxA/B7dyPBBymsqu+KW+8DaSiwiKEnxd4evFbYoTZVp
NOtQbkNu87y++cnJgY4FPDzNQqH/Io2LUQO0E8zl4XbKcLus2ImOCZJgb0LY0n7E
H+IV/t4FCzBBWZLCEcK1X4jfDKG2IZ//T3YrOgSXhDNEqbF+bcz4yiKeBMlys5Wx
FxX3qznfTia1OJC+8fbbm0rWrC/q8zQ1tacUO0F8wM04ln5vVt1Urjq7KGW5s6V/
nwt3qwRenCw3s5ortUDvF9GJGpt7I5axMAX3BkrK8AeEowZoyWBJ47ctv6li3yvi
6bI5XQPxrLdgutbwFQRKq44sofSvF5ZUT/mBWNgn3cdYTzhs2OXQvyBf7qgUg/2Q
IK1dbL+x3O6Gr6VacuPOWy9is0hgtL5JdsbzK6GTHHb7vmCAl7Wzwq6aif6R6NPV
6fNLoeHkRN9PkTOKDIDynnKKnzA56AitUSmuFBGRSlKrWbKcVlNkET3bEFP1OAtg
BztK02h/qYaDVbCsoyGRi1rpTYvX+KmRauOFxSsg9t3rwhyKejV6EMAag3vcwJz6
/yqPPHbhgBvRf+0vD2YH3MoNUcclNID8Crn7YyT/qWa+0pcPIz21yKz4ynZcQAUY
ZuPK+KwK/aBreS7lbvax+EYwphSgLWLVx0dsHgAWifcJSFdS3NT1fPgP4cmQGsOi
12fUlJBYOzF4L6nMVxiff3/cfhJvGk8V0TYpCLw+8TZ9bMdHpO4dWAbDHDIWRWV2
Rq2tNvUzyf0zPlDMZ6LRAhaE8s7408nwlYiJCdTo9HTXwnSNJTyJ04ug/NBeFWz4
/7GPcUFoiQ0rSD45S/U4quMu+050nWFnWDVbVvtAwRlvMONu+6FvCotxVzJS2rUp
eyefscnpiLOpLrZ2TKjXUtqeic0ksTn8KuH20+rjRpxlhU+fH5V4fAeQITS5yDym
zu8EidC849crRBoLm2TDkz/GuDaNIX4yJdCHu65OBtZGmp2KhFn27kPNfjhkc4GR
I1fARGEk3EVo8ETDyz47kDStl4sq5JjaqaQ6vB9RlH/Ce37wHLAePBjbUFMpzCzP
Bu2f3TnemaHpwdOkXNaq07iovhJzcjPyi+tiY8a8lrjjXdeykSlQ70/O453vZEVo
QfZ5c7iTT/uDht8nbvgU9JYHRTBPv+yYjtSFGY8yUDhb3RrWf/sTl4yBZzJrARtN
J0I4TjSIg7LT3cobQ67xr9iHOl29ymEQTrbSKXKR1ljOZNQmZXqTykhxe01UnNkC
UGafRaRY7esRg7k+KjU+j0cyVRh7GSxL9vqHYf5gv3dZMBE9z6w9O7QlkP1SW/zc
cbOcSkvshIId+7eQNiov9TbcFSlMGGWohXfWYaslgiY+6yUfjjCDgsyqdth+dcsI
q6ajpXdDeA9zKiAaeeuJ13FBqAjcuipdN5KqCRR7G7TVkVyJL/QfjFYIHgDyNUF4
LSs3tJfhDUWlSvttLffS/tqQUP0yQcil1kRowmkJDCWFVAIXhBeGhHYcqx49PKNQ
vbwrwDnCScT9jdJzqYmcJcPo68J1BKT3sAaiZADnPly0HgDk2w3MRiTljCthCcXr
sJSedNtc0GzmETInXtrAw/3jS/4Z9mUp+Cxw+jDfxsvYRO7hOm7np6Kx+gDAxPkD
6bbey5CyrIRYZqakTKt9IErEdW/wGzV1udFfeP29yUUKhvQc4E7ewzvJ7WvmvW5h
khz5jNfqVVf8FExnzVYnI8eIZrwnRwnwoM/7rHNjKH5dYyscfr37Oc8f7uXYcgB2
WSJdNfPqVpsssv/WNyhftlyn9bXSd5mHsgZm+cSroLGQCU5OQawfvWe0PYswyVOY
5YwSJa3Qbcw+QmafSamDWLTDChlj9+MyhZ6YnsWfMCGdp8lB/8KEpnUquoJGYF0W
9yFloQ4Y5sDyaNfuvPLOUZBuuGKYXJi7U/NLXSMaTF0UXlMr/IZctOkUBdddr3zg
xsARTqDop2noDBd4yhZrzAgFyFVNmuJsblQUbnXRsi794uEWwM2S4vOO1z3Lx3xP
GmAKpsNiQBJDXbZT/IH6w+SjTqkMMj4Mtgb4y787OhEjm+ji0c2a4KxE5S6J5T84
82Co/j3AfARZCgcpTcjYTqGZvIXCfQxnq73UoSIoxmpGzly37uEohUyK0iRfJjtb
si08Kj8TYiVzzctuMWPJNVJ83gtf1fefoWS5REAMKmtPAc9823F6APwSPUzlMWoE
q3MzpedWgVS0yMpuvbKwqtobn4T7hHJYTdZiTOJTN5X0qlz2R5n9BISGQxVptk5E
NCGwIjpZmGA2lisRmbEvKQTwZYyem4WNJbdWJLtTtmhYOtY+nuZ5KRZCGoiqY7KN
vlUuUN8owUAQ6gwbdpTfFZDv40zP1TCfqpEWbcP71LJ2JJ9akiR3wyOFwLBEnPW8
K4+5Y1LZepJG0lw0j7jVkI3Un3qVMtIHu6M+LzRIpa2uSeNj74irVRxWSEcDxDkX
kdDpZewnqrGx2B+0sIuyj3Oqei4j0rT3/Q3GRd9u4aCNlng+WAftpmst1zO7Iu0r
B5cdclzJ98JzCw9XSfA6owaOs3mjr75Ntvd+2be+QUtv8dFiU4Jib6pkaJaU7Vim
RxOj4QNGzkjsTeq1lqkaRyUPSLXn5gLJTTYEnd0Jh0CQ5eXB+lV8qOVMWPm1kO8n
QQ6+i20ZAfw301pn2dA7PR3Hn/q0XfIfMr18WpqTnNO3/ycApbDgvEwppG8uQ6js
wmVRnOlLC8rPbJDxEbCwh4IKefL8KaYBpJK1Nupm1Z7wE/Qm3TTKZaU4Ly8AIhdZ
L1foe0WNsiHJzWG18YbKQHWBNPXLoagMUnNNc377UjcjahWQmUKQDpTzB3PjXjBp
rv9uGaqapbG/ZrYDfLVAUOx5E0WmXG3G3xfTgy70p1/juGLohoJgxAAPQHJ+7GPE
eoXP6C044J2k8rVXc+2C29ZKYNqyTs/NxAu+OH29y7cg37WamLBeIenmHKJU/MQO
JrlIQgmg5/Jt4VhWYM+0Qb/o1MahzPcVZ0o1LsRUNCuVfnhydvGHLAKgSVkULFhd
x/OEdAIovDQNfjnYEtSXhFEDxzU3A3Tv5h6xDbrD0ajbfLHH74cmWminjcIQhOYh
Jsvz0S9uzCI892er/N4R1b0njt/OdmJNiBIOMGvFzwTj8+F5DpOuNMrC4JwCtHdV
8nakvzLolouKnLQbqIdwhbwFgfvpFXwZqftLhHi+j7pSmLrYJnLTC7Gk0Smh3+0D
CU0ZyM479BEDiRqodcpsD1sBerLsblWC6FKPRkeqG05edA33XGGvxT9+9uCd7snK
6SVwAFjwLcPtAtZC36aOaTaBt/VjuaVfEFzdRwyhmxKXsnnwnltC+jI391hlOORt
IzK5oFxqlI6YLY/hzPyP9GuifDnXy+87N/muNQPpNLKB4m0waUCJEk1JsKGYtWWW
we6W+fqS5NnncRua6938eTzeFZ8Oyjw/imdtBHn/pdvcNR73+tTzMFDDDZ9EE5mN
YMoeVYeOFgp2gaUY569QpQy92JJlsM5bMumPRQ9F1UiWbgAWemAyYsK6K2ZCQGnK
Uyd3UtnnRD/t8W1Yau2LS53bf6xHoTtQcjqJlwn8IXB+VcSFpsKzFGpst6YzCCof
MR1Pg2+FQTFOlv/9jhoiwWSN7qes6CWjBs0A0e9bsopFk1odiX2vMaq+332MO5/w
Crrj+SziXJ28BxfmNaAPXDep86uIR8j3Fe0OL+AO2TLNtB3fi/rbcklR2NBqjX8I
mgzfa9PuNwJnTPBXNF08SCC8xjra+Z8w1X+OezSWCTrPDnTh17BLYxL1SOk7aB0V
zxMZEDj1LRHrD8+7yDBDgbN8jMFghMhnCEd00OnCSCZ4C6AqXuc6zhrB/lWW+Dzv
QnsH2EO0UqZ2jyqPof0LC8WkZ0wn5hsFLtuT6bk5Un2Xy9pPikbcDCbszrwYpJia
0x2igURCIqHGM5n1UOQMXJUc5InkjcUluKUkXg8BNUSJZGft8xU4JkqGx0blZ/8o
IkGCSQS+dQu84fvlDZcIpgETo6JrKhe2GLvd9KLFij9A5TxVDjVeiF6wC4K84QP8
iykO+g1I3MPqrFW8Rli5hmxjcRwFEUpI6eYOpJmFWLEXQshJLa922rRAoerr8ZnM
LuKsorlXiJyuJ3es0MdRpp/+YEl473Pf9tX3kS03zKgv7coyPIGLqhMZdtvPymhK
jzBEvHANV/3CruRZc2T75gumMiGlFGuOjGl1u2Jju2geRdAXPuugX/6QGM9hikZN
bh9G5me0+3L5u4kZv8IH8atHNBdj+mtaT0/27X+X42s+kRrDn2gNE6TT2ZRZ9lQy
eRZ74J5n6m4p0OXXsfyv+W8gYI+dbD74Vcs8uB+2vycgp1M1M7pvSFnjVYPBoamM
cFfGPA4VL4WY+pskeY+2OEjfU4NT0xKHSx+bP9CQD2V8IIhg1nMLUnJtqPfcnNra
Nk1VHxdK7cIa9SKicvTam32xVgV9FW4bdo89M2Ll4Kio7nzHfPtzF9PX7jQJOaDI
SwVtC0ospi/gnYJq27L7DCQOup2R7FERSdynt/qsaK1ubmZivxAKA12ZoM0DZj0Z
S3eQUv8uaNGcZnujmczgsYJaTAkLweLmMvyMy/Z5qPzYnFdBbDI4oUjHFyX47XX7
rPAfcuBZtSlgbhTUihaOFevKGlKLB34cyXEeaKZ/DpQ9Y7bXO9swDhm8kknYm5Yk
nnmJtEEQe+rnxBYVP+Hur/9/4i/vsUCKlZF555aVtig6LXj1s0A2gM+ygZepF931
eBg7nZBgc+w/zWGgonMbaBy8XHmlHR3beMBD4PVDwbnGxDtB1V2rlkfWfKly3ePY
4PY/LtDDVHPdpN/Q6rXFiVc6WAp9Wjzpwm+wiTJ8EefKu9FSYFuCYDxKnifNBuMY
qNb8lhK5yZG9Do6eSQYZkLOAgSPLchjXDnYMprPXU/53I4b3/s6S00CzbBCvzQqm
yBwescqxSjzfJddKJC0miIJ2i93PZm3AtAPOBE7gt24+5Shk3RIT4H9AapcfwLKg
oqLGYD4rdLODMA2VcZiQa46tH20204zPUvrfUWgTcCyqEJKbqqjfydvRTamBnHHi
mMbYxcPzYHTcwx/87iUEdaOdZ8Be3TLH5Nkl4yv4g3hopv1fixQO8JfjZvOcA3fd
RoxHPFD1Rm2Y+TuS3Ey6IsJx6k5JRsjERO2t2cLL8faqe4emYZ5HbfodE3M3IORp
lJGWlKSo25/pcxKliaW/0Dt1JVf75ocO6+35MZcyEP3ZiOoo7fgRuz+dIv+fqwPJ
kuvH0m6maKwfH280TPxAD+yWwPr2IgofdsG0DpasqCFZq4Jlxl6vHyWShPxBw4Vw
EK4N6Ukv6UUlDodsvz8QikhFc9JmaTDGBG2Fw5vjlef/VWWdmgKGk195evSp6tjd
sJ9YRnEjOO5cOJjfjCTSJVY5dn1pmiaGeH32dl+sjzZubwV8KYDo1OF0MGTAGiOt
1aIq8GJhKnEMSLdx9/uxSYq9DIymZ+EZ2mt38iYpVWl8L7pd3cR0BmfgLC+tzr05
d4YqENMch2iq3IwFlTLyHdbaUCqKn+IL1/YjgRjPOy9WILPsRna/jyCp4hUEA64A
+aG2AtfWKI/I0Aq1ROd7FDI5Oxf00ozJM2/xElp/qnSewC5CluKLaEIHv8w/V+NK
4rhl4Gkwr+JzEmUR3BXTfWQPB3SdJPUShnz+Ot+C2jwtvdPO8DdKToBuQwIDUqM+
ypPyvoorTRDBx7zkRrrd8JEoNek+h0ImMju/dMmVNaW/RiISV1vweifMpOwpldXK
p7ZHruwsUa5sQAlPC5THY+eONQ5KuKPOEPjp6RzyRJXzn9v+DcJhsjurAEWWGQ4f
Cb5v7UcpcBjHz7bXZ6nNHKETlVgIbxSMcvTBYVtWIslHDL9/xIiAKxshyuc4WHqo
uKpsBQVpW6ZaDsks7Wl8Oh75m48arvb71gCfqloxZiHMER9AEj+Kg/9yZUtTE3Xu
1vHWmzJXf6U7FcK/OpxKryuqdl5SfThB5QYQfIS0yfFswaYfPzZyV9oteKuXpOa1
btffSzhWVhfKpr9BU+/fEsrmLLtmpIeJfLIHaGlOL1zoRWtmM1kEBuTPUi7fbVBW
SQrIDepgRaXUpSYA6tvBJFA/U1GnkHx73NZt/rykK3INZb9WjfXqeAM+fsLc+zAH
aIZkaJdb4tvDgVFKY81OWAx4VF3rLDw6IwQUDfDywgqkuM+QFscJVUMmolqW06Xb
HTXzqETqfOIz++6Q2zJ5clZLB/PPbM/bY1akM9jW+hh8cZIJh1KYYa4KIwFNiDSI
2APmNQQfM+nPkYSTRSYzw5H9DUudceqfTt0g4VdSbVB2y5BUZG4cZ/fpcw1LiR0w
Bs7wUg5jrbsCnnjnRJWrPFj4v7MDi75yI2AXsI8oga/0BnDakApPIjXGKU5vah4o
sDWXtMXSFEkEiOVsqcGAeogQLZo2YIl50kBdsVRMY8nt6zd75wMyjbE0z7Ogvxvq
LBJBNKJNpIEznLwDFhdppa8P+IVHEg9G4wxYvTUFLo/L6UsBF9k0U9dLd2riYQC8
8CbcwcgNNlUffPkDioQXtMAbpOcRYK+l4c2mRispRJ01FcGbvc8rsvzobEV1V/J+
WH7rCRI5jHq1Lhal2r4gl10oH5wI4qoZbb4vZQYh+BPBXlAbwz8mbZVmPKX9KKbo
rk4sfAJtyRYCO8vPpl586h6sOL7WwwmQY+BHGSAQm0e+0byevDuhhR6qX5cwdreX
HWfsQUO1/TWUt0PdurFIsls7RNy+2v8bsnUqTPriL57kvH2S4Xf682tOD2RnLJ90
L6ri5wGBu3MgC7GW8Q8Xu9NA/rWyfWfRiaUmQ/+zc1u5E4DxcDi+XGPYDnKrHP1F
hCKzOVcqJmUc65w5q19T80HuEY3SlkX0Ybf8iLi+ASFjdqoBnErbg8AcAC8GoSCz
YcKDBHYi3weNRxsQw9lUEjtF51eth/EX/W792D/mvIUhQnicR0p2DncaSEuI7Wry
8OedyGNK3I/FpINszQpJ+9027RDoLmd+DJRk/pPqfX3aHp1yfajNyOJ8i2FTLlIr
VAndriy5Eme8J2rcQ/+qK8nW4i872Sreo12ek0K9PupHzDc91JRs4tw7d2v564wb
+1k7HSMe1CGSXECuSxzWhy+9cJ3kQiz5+uezrnqzRCVBbwYZxF8IVfFYZKGVFU1H
OlWJS0ftIy3lvIVgIeHcKlA/lAIyFpqCSiMG+XDl8qfw8lOJfEZcImHHDfuaHMtR
lq5b0J62CsW9fELAbbsK8cuLRw7tKjQJmQBXBtg9vU9jkT+BKYXMqeNtDHTgGyZf
L2YuAGNJklA08TNp/Sze+RCnHIQ9Eipa3jkoGuDsaE6Nmzd8VFkz++jBJG5pkzPA
g0340wsOYthep1bV0gz8mvsymuRrP3RgsHzxH+5RdylqRXEPpsCCcgWg14D2xid/
nf5G/n8rp0dEjtybR7ynbynzsLPKq1FDqplYLMAULMaY7/WVflM+RdP6mL4PW2Qv
3+OX6R936NKA+9L5pUrqs978ZYCS9L0pZz885pAbELKZ73zqHaFOKT17WP6q3aSm
hrf7Nm46nmwJRh9C47ZXPfHBqqF4duHNWxBYrPWlvu16zcfK4WNZDAzZZJ7kAKAR
9UV0goGv8+2VxpZj77B0yOTxdtrRzD7UF24pMYmqLl9qwESuOSFEEqyXfyA5neNQ
eTJHk8MK+cslvt+lrvjp5RST9YKeLuslBw/iJydoPEBWZtjxcH+MrqnJR3q2/fda
4R0JwiDWZZtnSxcOotZKR/nsLrQoKOVBSm/3kH/Uv3NKH+UVWKYwzEiEyEfVWi7a
NosTZxX5xPN2L9ht++nllFlaurM39/bFf9mCFB0TAsGOJuE7juTWnozlwG5BKh2z
Xu91+rMO8peQ/hDqnQEEm3W3J5zS3O3QM7JSV0ItSMRcDKyovAdh/UmsyYCvnRnI
dG+aymQaAofSNZWlB7zq79DYzDQDEPxXtg6TqOgT41Iwt6T51iqTdqlIt0m6Km2f
XAwNd1O8NkiZfSDZlTB59NtggS77ZMekvSMhGFNCfniykofURg6WCFxig2XfZ/me
dBQgNz1MBO/vMpW8Mw/ExJsjA/pvZxH9UaeQgekcVk7ImSDncVyc4UbydSpiKG4R
NkQgX+UfIhcEmi+ZC7NglYZRlW2CoaaDjEzzhIrBXMrOjjT3FVqJv3KJqJnKTCuO
UNvVXmWKFGxwvn2eXJKbG50y8zee9h2NJsZZo3OPhJ+Gm3BNGqatAdm5uNWWPcOp
xPcuGhydggxtkoQV0unT3HNLtpP/HVZtrL1/qtbD8+M6y+tsT2J9oQXgUxKV6YFy
KdDy+cci3Pg9bqi6UfxN9aoQaNst0RQRcNS09PHCRW4PC3KGZ4qGv3ykopovcSRV
ZRx5AFIlXBX5vDaf/akrRibphkwKhTcmOOXNR+yYgys8QGRE+85k6BbMkm8jt4Dj
g2j4C9PusSLhU8R2igpa8JX+UgbbhMrTAfY2V6S3xP2wgOhduzU7IG78ZlNGaZ++
8WqzAU3GkqNWmvG2AxWIxcHRPnRsJ2SEsBpdQ8RrZ4+9rdTnrHF534SgaYO25MtK
OgAs2nkw7pfBhonMji5rKy8SMqUarwAecGpo/OEokpDOKY5TiA+qRhCGyFRJddbI
N1nXZg7QL2nPtu91IHrXE8EIY+0bOdli3aBiEW5NKwu+d9NXQfIPTNJQy4/i0pSM
rzwzEICq10hoIDakZL+h4aajbOgBFLRgjjpRkrAOfUjTRd1eUUXgtpIfl6aJBdDy
7qIA66uf8tlJcbqGqubbksta1WrGiSBtXRCHUWY7qYXmAjbnSfhcQ1MeMXZ5kCmf
0NDiXcBMbJQV7wBznnY0x9I4jDfI3YuUzxpPh6+zE8EoMO13Vj/zoNzAIIqreZr8
nSKRXoPGjuP2r27Bi5Iv5aSyCQPm72SF93jLw42YtrI3Jjd+v4wF8IFmHRVn3cYp
9OJX3hZIp4XGQ9jtFnNfG+M5Za//wldDTef38PMiT3lZJpFGYtPsWlbtt3t0i+ZK
Puewsn1qq0iSsGn1R2l/wGVmVMNhTahUa9JdeePxlkSXrRkU0LctUfHm1j8xknHm
H6+P+intd+FbiGNftf50ARcHp/zpSSxOFCOF9ZG/2CLw29v57eifUiYnS1Hdhnbj
uh4BsfcNPhnoa776DPuO6TA85K6H8KklQnrFbGYFKCN+6iNJZj7kvamUarb6qgd1
HanKUg/l3M7ofNlmtkBSChxo8TRuFSoVI7TyyS/5S9xIsAZfdDHK3f4br6an3MbI
yZem6gRNhOtyob6YbNEmKd0x/C8xWHvQOUqeISz5GzDun39iQTm7FNAYiXrGdDLp
VwK5bEoKUPSFifbiHqIcT2tQPc/XIijT1dL4qDeKF/6CtRP1biJhkHpSCUzySoKl
DYwWWeqkcnIhVj2ANkaT1o0Sj2foNb0FKinbtyf39csq9dSM14h5o5ecXy46Hqmj
lnB3jG/ZKqZbt3t7EGk/qr91YQzVjTAhsDll2KC3qjeRuG+4DPZp9omT2s2AdF+2
Qh8yOvsfsSstol+f+ezupJf7sOPVqT82wDZ4OVFBnsZ1ykVIUN7KtQLlTfQ7bRsx
ENfIxLAldjPhHZfUobJESZ3bXbP1LcKMEuhAh/5MZndQaU0Zonb6XVPvzteG+0o3
wT2eRbHS1+rQ0CpVKO7IyVFstQVRoUQtW5UOY55zbJjgtDkuBVcl774ZGymv2lMN
ow25tkc8C8rkdqk1rqyhkUayqLAd9okh7lDuUNJKlGVIU8SqyRee3Xb60Og0Ms7r
3EcFvHSipcARUlyABVA30HjHo4l0aJlrzNmD4DtuT1YkIFDe3nvutrzmUsH+RcNh
Vd+3HWxbV3dUAIZZpj8yHZ/Wpt0zdyI/IuWZBxL1rrPVRoerBhxwYdykgoVNoAK/
TiLe4Gy84vXDUA8jWK56WbhfrHNNk3k99XA1mOZiWIau8a06+ua/tGoDdDrqKzwH
BUEs6nqRQvNQVhioM4qtoHFnLk8j5HRzwbSJve1XBvhYwdP4ST1rOMY2NJL14kAT
nX37SpVgLdEaPqtWxzh2QhennQjNEtPU9QCots1cCTuLxjbfkxxz++bm4ClkTWpa
TgAFb3xVrwYgFsxSYJ4CZj3toCKC6SurLW4jYiBTggbSvfRaW3s8UCKUEHUbQV/y
dv6RbbpZKGKmiGzycOgiWgCP2ixh2aiXAnRKMPJiWwWmykp1FaRdDO7JSHRHj6rT
TvYppL8N4zaJC3yd86wLojL9SD35DckmGO3Lx9yXBSGNpPmVH7GgvKjCFN1YXnj7
tJ3hD5quylnGwA5VzytWBj6CW/nL17wrJgcALPnXet2KQCxCi1bjDXje5OQsWxAq
8KlAsagX0EsYolBePbb++pDT1W9f/56NJbFS8Xrfq5cKiEQUdd9GyRugSPAoZI/z
PWYz6XhwHrrxzU7zkni5pqH1AUqixkJthyh6UObYQ5lPRJQ51t7zjglBsDQrxMej
qIBlC+Sgl738IimGexbm2Y8qJlf5ZtecU3mRY84dM7e0a8SezPsvnF6BY0Qy4hPn
8nHMTLnoMpo5jrajD7DGP4bFhuvxYw4l99GntES96Vg8fgaChlciSYncNr8mhOMf
MZ+dGL7ypLv1svZGcY0TGmPU4z6JL0ldOssRy8qksh0Xo//WD4IpooK9gZI763Tp
GpEZVIqRczFVq8qWf3SbrDy4qKsW54DkdxVZDSTf14HPv9DKkKmF5d/Cy1BzE865
J5PR1DDQq44Rw3NWL6/fLSIxmgN+m19gcSrR/Xe8UbRB/p1E0ReDFQ4dXlooMeKy
uXGRvJ4YWNoR9Aq3I0iHJEYJKXQ82Mh8XdHd0BGH1tp7FhgXXR+Z9k4EsiBAmhbS
J9/RohECbKzWpgBnxC/cTeDIbwq1BD0rl3akY7SruoRSuJpEiedTMDt4IRbamg3B
UEE+MhBd45JLVIA9feKUP68O27odEPhseA30Ss6i+aUxaxPzAhDB8U1g1r0ITCV2
p+C2UzpHU/y6KhNjiuj9sIVCffTSMVZxCtn3Ub2cmMcHtJiasBFcAzI2XDwWbvjZ
sJdotbK14XoxnDkqgJ6wX7+VJikAsMSKWJAvxLgTKeZyA61byzoRaHRSw+TasCiI
0IU4Qg2ZkTfEoUVSmtUZJKyqiAl5tBSeRbkgJWcUOPxYZZ+wfZrV8rylZElhS2pj
1LdLAfevcoLx+dB/J2HFAy+RJWqM2znZ7Y9a3N2vpjGh+1VyP6yEFFNHX/mC9UIu
s5e2C1blnuhNQMkxsvECbdHhSWkDe2cYB5gb9HAoBR0mSAZEVcPCA3Ilpq4mbrsv
KobQ8xWz8UTb/a0gT0cIw43Q8hsiH6QuW1It7+/C8Fc0OAcp2IKmtb/JT2gmB2hi
Vp+ZHvF+3SjhiWGSvLgBfCeAIGPHgm2MbgZj2yjJQXaI5bGn6ZaAO/wc7cmGC6to
I42bSVn0/KMMxBtyDMUDvklpRBMzvFtT3FZRBVNtasgWgdLQq8ssCWOZgXxQQjPo
H6Du/GSgr+8ivZOv0o4wc3LqZDT+2AZ0ZLEro6bh8B7FaskqVCKkGPHPmzz1cQxV
rlAqqMAXDxsAYCenzl0TmfS4HYLTrQ6XcQEFyWXXTNkXwBvazr2zuN4hGzBTLVqe
688EhBAS6RZu0tp1Jv5DzZtN8o59aG2o3X7d+sXO+AhKK3vNi08dQ7bie0vTEMqh
TxUmGTsh2SRhM+pfUtZWaDt6lWh9xPOI0t6TMbZwzIG+vnSdGld3LO071pxjmrxT
fhTOJvBofsCD6uXtyefg8NdjTPOyMbbGDGlSw2MzUaSThTK+8wT4KMgp3fdJbSBm
+bpv2qOe2Xu+VO3jt5bEU1C1rfUePsKVmjth6GsERBfgRAL+/hQcwWX1vTb+2t3S
q4QbSOb6RZO6Qx9Vpd12otvYmxWuglOYPtRsX1lpUaVzN5oXkf7uyIUJEKgM26jW
1pnyZUiw5EfGwziW9oXL3zmhuPaBRJStkcdHJHVtXeEJlOXqGEeXYmHMDJX70YdV
ij5y4qztC1H+PlbCYD97Kw0cVuy8PwZmImYIsqX1W126PFZfv3RdZLZJ5OujduY2
dlKnKqtiyh4tCUhghMlLUsDD5jh3YHDate1IQLSwi7y7/GAeBGj+9a/7zDwTnam8
cE7cWcXEH5dibJCb9NrXb9m1JpMYHinKbCjp3Clj7mOENOWe7owcRj7H2rr/FxnV
7lnbDqhLPZ5DFgc9+lJwOVRlWVOdy1zF8BlyvNyuC/PZgnoP1ehk9871sLD9EbzS
hk88aVGmiSu5J3qLFWOuYTe8dLmOC+WTa9Fc8zSJ5xZcoXSpCBO5qY44IWuQs1Kn
BntH+j0e76BBMWXmMCZQaUQtrITS0b4DBc+cLB7/Mga9Ktg+vxtrsiWJr1ZhFfbK
3dVwwd2G+JZOBqYy2um1oFlcuFLmQIkoHC4upa/bVWOhwzo3kTKErHBTXMD/Fze0
Z0h6n0ayJxp6Y9tnJRpCqx9Oqum1uNUXyHKIwAt/bzmgBz/q8UPCTzYfoeOerLwH
s5axIFxZBkuEhHHyAb2vJWiMMm2N80mbYbxaWzYo3w1rTc6B8h0+3Lbj1shMYqRx
zZlg4AraKo+ppGe0wPbZdEsuLWuhkchGkEk9aOly6w3mmXYlH+9wn9oI1ZyS1yOs
dbACZ+oGHvoJGpmlsLFrf+al5kji9bfDD9OSuq4q8VyIdNswJdwpKsQIc39/T6m4
33x/wryHi9omib60fYk5tHk+DaGdNLEzcspQpyyYheqgq9jfMvtU9tXUuugLLGdA
qVRPcE5vpqGN203+ENyZDIfj/vpIEPaU6u7Jd99eUp1VN8tpo+FuN69uslc2Qlzi
uIFYd0xPyyMDRWz4MqNecXLddJur2oQsdvTynOwL1iEa3C+/uJOMgdTGi8MZYmwW
CRV6QoJ5SkTtdjI5hmbmIGBy9vmTSdX8jl9yZ/aqIEiqB+PD7ZihiKc3ccNiEGdb
AjSO55enHfZLp+WiRFbRmUN5m1TI0zqM9a5ynKPgRgVi7/BXSHXGtix+j6xCpA+l
XB57b+Po3/5+2Hy3m559KBOxXJ+lFYUkYP1ZHavpeJPhOAfgYTqySaO4ve6m9KZd
X5/JSmSXU45HfH0U3c+QH6VefRYpNu9nM7E6FpSWM/a8DImpThqyTEY7AsxYjjCn
7tS6zsfOzQioyXbk9rse5nXpOdcy14mabCirwvC8Q9vqobpF0hKHyUu6WCdcNw0y
Is5xWB/Fwn0HubIxkpn5qhlS4vQ1GJzZz7r0YiSjJ+7eE0QImE9a08Z3/ZqVhAbq
kXgBm907VZznz1OC+D9vkr2PORhnDJ87S8KoofU11wqUYp4x5LlLAcizKZFDKsVa
+BFsc4pnR2NkyneCIJKbRnvsZejJxTJIeA2zl+DovOJ2dGeocv7Ag8zW6vkZKLTl
qdz0gQI6GjDOtMK3/bSX4MArYUUE9Og+pAguxrqGR7dVNWr1DUPart7+HHMgz22e
ANxGD7SGz4jwic8nUPOOJ4HRRvhmncXZ6J8ogrPT+SYOjiUJIQanQ5gMpcWa3pEq
Z22r5Wt8ZQGRHJJBk9g+KMXAgM6D+hxSmTag7kLxm2fl6yHffgR6s2/+5LlXGyDB
X2ECBd1OrMBJoKGtCj/acnSL9k5I6bkgZe17/9S+xqDbs+21p0k81AwLMU1BP9Bv
r8sqz+HfyAVNAFuAiI9fnMt5QJDyJ/S5WNVm/E7PI1Jfkxy2UQU2fs9wzrmnmpUU
HU+Tp1qGjVweoldQDD8+nBr3LnVRpoZ0hqCoiQDT6K93WHnmVAsV+IWkSaeOtm76
l5IrDU60Lh+8m9jLN5312sfJmbGN9rvRJ1oILsWafja9pVjUtD5xFv3D8kccq+4C
afoWOPrS+eo4MDfJvli3K6xe2CmUPfDiJOLFE25IpSZtkKggw5IoiONVOGk5h/4X
vqqMgyQ8x4zZugVH3pNkuU3sdIfoBsRHurjomikdMgvlft8UIGr+i7FmJ4hmoN7h
xQ3I+j7+jdIqYEVHn26+N/o/+/xg+q0uo/P0w9Ei/DhyCEHXf+sEq5/Lxei13LCB
xZM8fvFvYSoDdkZdatqQ3ZUNGyMFa6vmUK/CxYTiAObHerOOd374rplgOHc6c9lV
9/EhNOZ0/eYLEY0ZCtPnli7JCHDHo1x6PqggI+fugTrKG8fNgbucV1ffH+u6TB01
6U0JsHnRt9HK68lj1mQlGVzVsI57tyiDl+jc8qyjWdgDQmOJPeip/+b1wYPCP0BM
739tqS5470VCb/HQkzpeVBOscLLEIS+BeuYnjRJYY708Bvo6V4OoSovoQy1JQTok
wzyVcdpdaMmdX5QFUMp6sdYYXHsv3Sh0ZWylaVx4CJs7PJIWtBb9De1Q/uJnWtc0
BsZQn3b5LKdgao2j+zlGi0c0tNxkYOgMuG9NIl+ZElqxO39fxc36YxUlgECNheqc
bbfId9CvIGE6wlGSYI8fSw6qODFCJMoBT6XZclr+cnZ2/FHaZVd8/NGgV9jUxrAO
pWX9BIFeEN0K/ru+jOuZ7wgdPIoCVTgEM/G8EzVkJv2E1p4De+OtREF6rWFks96m
5MRH9Jj9dJWoj9ZwUNpULk4/4WgCP5nlGVb+Xgo7TscegIDD0AUDJ3dsOiMu4bQF
92/j02OH1SuYxu0bLuxvmDdqywU2KlJnnwrMwUx5N7p8OzDU3nP/hE6tlTYIHD8K
ys1SZSGjFsQ4ec8iYTG8kr/toVeQKxlF0JdSOP8ss8la6AJAUq0OE9Pp57mWjZ/H
nSeiU557lgY+wF92OZubA8xWuhA1kR7bMaP9Y6ge7sFQExJI6aEZ46rIMczu+IEE
okbuaTxS7O+8qpq7364hIe2b1Wrm6oDD8Vyv+dbEFVca1a9eCeSS6sWnnGOx6sn9
Nl83WSfI8paoxcG7KIq2mL+5YaeT7KOjCNwFssYygxKnapTDNli/HQ8dD6K4kEPu
FnvSCb5VCuYDB77NvwEGha4xMcoXARD+LalF7DebjpKoy3r+qbCk3+XEUyvtlwKR
ebKHEdiGRgAmp/NvYEBqY+phcMu6K7vVNF2QFOF5ea7UiaO4jvJ3Bn7ARnPHphn6
okfq1b5a5GeUQy3RmGynTJPjkMFqMb3GxhaCMv+vbQoEwFhXDxTN3fZbxhwUYMVD
KRUoeoIad4S680Ull/kg8z5kcANpqsZJhZohcbFzlU7oDgCOvP1rljUIx+t2l4Zu
+0bRDLx7x2X6m1aP8NUbhT5RUOEYPCNIeseWMCKLS2EkwBhyBnMRV7nVdYG+jGo0
dTG8UPr4JvP453SB2RqMZtuX6h+LSbGrzRl6E2hzN0H6VIoDwvaZ4RH2NVw4ALRc
JQ5YCReKsuO0srX3sIPaiJjjV4x2/YHF1FqmZyVpm+W2C/GDT8lxDun1X2ab7gkQ
II5KL4kXgASpQ5TODCApytqziK/1XN3oVBOU8xkTAT6f6UIs5MuDcZzZgbe+waXq
YOGhA8Cb6aHxmg01BCpLV14ZJDGxcKJElWyWuBIKe0/haEO9ezkAh+XlJfTyBInY
awMV/Nw6+rYHrmZReDc7/np3vJE3WvypUsXpZVy6opVRWwI0UM4vVtv4SRsyadho
f43xh5TIJFFXYKU0exi0LZeeU8uGPKCCr62bZYan0YxYxAyo5OgRYHmd3sqsPPUA
sk9yh0X8tVH4hTsiLrLjDn1lnL4oaG+7btOy5wwA7A5kzOlPILCA+hQFdyStam9R
yDrrxb0BjqdOaMdOh4YEYHRydTWVF34UQfoLTF+P6r1pDUytyS9u0hgSTo0Lkv/v
DOwDaXz23TnTfGtD+0SWlEMFWI1aLseVuTYklcaUSQEWTFEnv/P3mNeeUdr30wUw
0vpSY64iYdcjAoqTPWmfp/+QlqBWOVq54fky/ZwO8w0DOik8LRlkKqvi/wdP/AEO
Vwu/qQZ/sxzRGHXvXk1FztyeBj4+ZsScduUP341g7k8/tT7+HudOm/UhZrX7k0mf
RfyN5Y2s8yiVniLxPSO3NtcPiX3ttV9lThZ6F+gTeG1oWdvxdQfC3u4hyScFFv7H
McJdPq65uebkb8sT+ElCgBz25buOZxbYilYbqcjWHDMEjp+wXTB3E4geeu2AshXy
/ELSG6J5AQCkSabRBNkjRU8i+X8FAh8KwLSrSZ9jTwidoYPHHWKkoFkF4LmvxSeX
TWWe3yqiFYovYlIcJnxMchL/a+vxGb4FzOFfauxRZWVfeI4EfRzRxup2Mo3SROXq
b/cQx+TmB6vQ4ZB9oY0IRLLKmgBwpF1iYlrAeSNf3tczOKpQdxSsKMzFFmN0+Fw+
OjDv1BUxGjYBWQJ7+1Uj0mpibyb78yNDJCZVG45M4ulvNaFjgPwsOWBbCMcI527a
hp27078FGifweq6EYRk/emCthh/nw+qOTFpVZBniZmTek0aQK4osg2l6fPlxsHyv
YD1ISU7S0dLS/kFOBFmpaqSqKbMf7ofdztdymqf02jVP8oxCOdLpg9wBR8hnkEnO
IkzGCIEPhM6W3ON6YZml7hqBT246eKwwzet9agQoeKRNZqnyZvK1r6tMscxGG+Tk
7FLgdudNivYNqHTiHZUPvh70ie8JEfbOPjxPyLB48P5jJF8Swg1i4clhL+ZRLooo
ifqGCu73JUd4zHUqAqRifNTXcrVJ+P6n8UHT936ibgW4laXsmHLcIYNG9JmwhUCf
RZQjpD6YXhakpTqDKbJYQfTp/koCj9qsmyzQE1qAjbID7ndzK0pODtJFRH6/OkpY
69v/4qs7wJyL5OgyQ4z1Mzrz+FesPCJlHLEZ4GS3IxS8cphiQb2yJAWzEf4XVg6G
Vro+WBncXAtULnL16zcGJyGDXd3saCrQ5/L09ktiRv+acLLtFjqXtet9hzgMQikl
FZBkaOYnx+l2g28kQPmb72MGcOjiMOgkZDCY2rRlmug4HJru83+uOJdWdghmjoE/
7yeqU4T5i0gBsCHCVLgAfRlSAdxaCMAp/jI7lLDRfmRBFWhw7iNF5GxEqyC+VXmb
OLhWRXjlBaLAPY7g69IJ0sqB7q8ugBc0Xpa44aKQwRVLKM9vo22bdpdqUT3jJQok
xCvtAtKg8uQ4nNJPwiQ+8jGAplFNKAievpqAC0vg3wdsmn8YNSr3vWUHFSwINmWs
g6hSOcbyXBZLeexNrXutSkoz+Z5gxlUiiYzs0PLSgdnO3evo/qxJWcq/RZw4lem7
MEdbDqRd53M/unqomCLvTJZs8GZP04bESGUDTx44EBwVWPQjPyW99sn9dI1FxGnm
jBeXe2nXdf6YtTADdW/eqN8q24K3fSu8oZ1dNgqcnqCp/ElVJThw4Sqsz2AC1LXz
icsqkck45r+Vxqu8Av3J9iOWLlOHIKHGV2/OdCO9jq9Yp8iqlfECkbdwgFjvFisM
AaRYjlggBll+IOi+kuACm8EyM+C1VzWy/c+4ww04b1qTFDg8mMkpNY3XTwTnmSnn
QI+wtbNtezL5Dsm2IPxhOOVBQs+rsFraknHdlt6JZO+ZeQFaMGyCGObnJVEgEcqY
JPJFI8AdhBNzScMYUpFcYThVMda6a25zK5ziX8tZiBcJ5RYLGBjrjGZrlMcQQnzd
EBhZ6OuJhvuxVt33RSX8IYgi3CmtEkHnJKa1t7hpNK8K0Q7cWbWUfwiNxIJ9ynZY
l6RacYJXBoZeZg0aJN+GGqRZpw2d6bkWAmGsgbgzg+Nf4+bmsmaOyN+LQ6O/FSxV
6rXQTm+eL8QaJxa0SMocvRoShx/ReuwOljWnYkMN8sAL0PgYEmHYwnGBMgBS4aeh
JQYG+kjOyGG5GGK1dYO81syZQDEDuHksylMPS+jmj2RE7Qt55WlxVhMwE+qh3gHq
hXB4hz9XqtIqSuDkkRHJ4ZvudkSbbgDJ1EbM8pQtWsOBnupMEir8ySj+Mh/9Ijlj
7YynYTkDfOe8CjnsQQguvymShJ9b2jxKh2QAY5PfC3S/eRQrl0uC2t34gwEKnCv8
WUwd0aAP7dVYBg6+0Kgwo7fI9bv82BO+SVw1qus37wT1z8zC/i1Y3QiwjkQbzqUi
SvLwkwxqqFjlja7v4e5NH+0yjzzT0omVTe8tKszliInvjuNRZrNL0vNJK1t2+0AC
wuRKNHxwR8dc1v0jO3qviaji50fi69MXRJeNitv6UcLHbf8A84f0vmIEXYEbW77x
sIEvEbEVfe56F1YkabV5z00rl7/BTp/LjA9RrpLlzZHzfeRpZO9dwoa1qTABb15M
m25HfzzrJRZaJiRS2c3M/IWbX6KtUFIACXHT/BeqeZ2mr9yFGf9KT/CbFA11XpIE
FdpuVGBN1rKC1P6jFjRCnKKUmit0/Qy8KOLer1sSCAbJHCWQ7wGKrIxK2tr9cktk
nByTCFHoI+XiFBeKt0vzTVklHjOCbH8YyPmI9g0cuMOhT7D68e3TuzzL9RrHGi27
KCu6f8RfZZmX4jhsjc2KHQ3FJ99sxI8tSJr2e3Z0r6PezuEdZjvTgYQ0CTA1ff7o
+5kQO6FIkReyL8l4WGQ6581PlfZDwbuQ++NP5lEhh9rbdqH0z/UoWsq7HOhzHjwt
JKjjnHW203sghChjLAqa5zq9WhyzvgGGtFGOFag0DFdcdNaBdBZvllPQa5A/V5i3
Ux51EpuNC8YSJh6rdMHa42k+uKQmE60z3Mtl2q9cAKbO6AKCCK4dkENcVJ7NI45t
nR96htGWoC7xznzi3FDApLstRJPIZHyjuW5cqNvHydz17MZNUUkqS0y0S3npgx7k
VYt2bvmcdqnG74m4htg6hspnanbBYGwsoDhVIaNXxNlo4InjYg04+4QvPPQnkqSD
Y/GTd0lt903nRvMEk98feXeQ4EG6lfZCdcwoa+LUtTlwosYA1hFYqVWx6wZBklJt
LYiYUqiNBBHmdsXuJFndFuEpAP/REekwl+Jr3rp+OIzjCo6o0X6NaXuNeEnYfuwy
mMNcDO544nslHj2N8oekxIUdaVaJUsb/B2FfQwlaYzYHDEKPRTbVMNXW9NUCZmVu
Ts50yQnEBIPxqVN4JTbjTx1NTEl8cDpAvFdz6FEOgeYRcG09j1zaFVMk2DnHvudZ
L71RPw90ZW670avL2Z5OHN5KsltF9pAUNOQsg//cDw1btHh1C80NL0MGprP52ppB
Ke2VnBS/a6Ezv3JNjPNkvtjvwrXU6C2Uya+AfhwN13+lGazfCOQq3Hms2ZnPHtxz
u4zyJYqQTL78Pogx+lvAZH5HfF01TOcp10+gNswF8pUgl7YwtT5EUb2A8h7p2hEv
nT4jQFlXOfYLFytH462TRKwgLbr/yPQfvaKnJV8goM8zmL3AJLVQI9liOdA9TjOx
+7wEBmmg/OecUHcwUXR2Tj+mIBzuXuhfdRpmSh5rQBxq5MDJQqc/QFCzBmgva09G
pUt/Dv+W9pJmEwNYJu8xU3eEC/bIF7WiWg4Ar6PPmJmmaR+s/Dbaf7Z2r5MBel7n
f77iHp9d0diKggfZLhXOr0gHcvV+Jv0l/AfheAp6PoHHnmeTG9F2qqd6YA1BrK+6
nAzf9nI6PpzwCaWCbdcM5GYx3Zl/Vb2zsDkmccP+Zoi0vtLZA77turXZiU4PPMaA
Bnh4r6kucX8xUdTPv+zHry2+6vILbMAUIZXBKHZ197wzpIaUTsFTVwasC3mYANZR
EU0od4cqoYcj2Hn9tYGnq//hTQw7ab2FB/nlslIqWZ+l6J+pD5Pf84iTviJ9F7Y1
nA4cKAeo4s50dVYWS4cnUQ==
//pragma protect end_data_block
//pragma protect digest_block
1FYJyYuWe3iH+HgeQGaAUfJhZ6w=
//pragma protect end_digest_block
//pragma protect end_protected
