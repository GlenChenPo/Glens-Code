//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+I9iwQ232o9jghPw+plbR5tVA3gtKZE7KZxfO0EyeeUP/hQpP+5nLeDac6SdOi6V
i+a5d8mY8hrhHVkov7gYzgmUyCRRCZDU2eH2MIyjUDX02bSi3UaZmDKGjIAgbYVb
nQYGWqTxeAT5eaDqs+755oxTk1JlAfuDbmSzqT7sdQ4tbYne1nT8vQ==
//pragma protect end_key_block
//pragma protect digest_block
iWoTk2HeXqrEgOdbq9hLtsYbXxE=
//pragma protect end_digest_block
//pragma protect data_block
sCmra7auSyfwxV9hrHG1uG6hsoKQqTo1W4SVCSA/DYKcbAJ9SgsCChUa1pkefyLJ
YJaVlX2Izu8yDP4UCNh/iZk7BGpFDighpIbRLGXvcocIxs721h1rtH7eDPMJrDAy
f25H5+Hll3jYiHWlgs10c+Zb/cED7b/yerIlhtO2en2wC5i1XBy/IlinsA9dnE/g
MwyskQEPsZTk3QNSoVcSq0fm9z19cLzAWPaedlwEqNjKiURE6iWPw3EHLBNnxloB
Vmk6xHn59FvzNP2caQJ5gA+9YhzuqsqutZEr0D7mVROxh4Wo0Zw+Fm0952ieaG2p
bpPImcnPtiuBmDFobWgQ9XjEw+Puzl5V3o5K6HOpX2VPC4ajDI8xzwTz+EDomjau
yJoGiRg9J1gRvePVTbz7p5M+D/joNq2yb3bIss7WXRF/pl17eFN0+n0TeDPjKOPJ
z2mpLgkmTUrVaE2nWF0+aJrr7kozp5QyfgJgm/mzp6FfyX6Lf2PDjnmQvXkq8Ma1
UFRDVmlQ9yiwlBlGw6nlMZ9Vg5y5qimcJ37QwhI0yqSIrSXU8ejYP0odNonejVnt
5Bmc80ADF/lK1Ko8PdEIoIUkMnCYh4d+9EdCfxIDqaXRFZNKQsGN5fDacx7nzid/
HUjTYvZMmDHCY4tjWi4gGbv+nGK/YfkmBN/5Nzq6TeGDyGsw5oJldbN0Z8Id1gGM
7s/ZlaqPPSNImDiYd+39AGrkKpOsSFpUbfPcZ0MzwthW5ILEcy30Pv6ej2AsmtCR
Ys84WOMNd7SaEWQP9vNS+gnes5BYUkNu5P2nDPXa/pYxgUQzJcWpJg/zXTassk+f
qC3Vf4y8Wk8XSEDWICAgdDiVrudtBxlRmgkI6+m7q/HOjFL3I8+ixhme8NIF4lxc
sAv/fylU/MmCC5m6/qSuNz0iCxFeYnzSyuyDSDqo5ud7cDnq5YD993MT762FEcbV
KK4M97jlGc2M8dY1f+JjCXa9sGitqAoquIGtD+irih7XNnmCSKqqJNI2+dh9wgVj
W2n7CembZoLSIQAaVFtEmZB4vae1lGq/OMzNkbci4XW+Jsn0hcy/n2n2BHlHNxqD
ffRbNSH3UBsucGJ/b1mjp3IMpByuLOF8RmjINHgTmEDxvVaotR/MdGBs2vyrW8eB
Gwwu7r7N/BUlftZeFFIGM8j+7dyIOtxfCTg2QwNJIr0EKzqzZ8ZiwnRjiNwVkT2o
AzuJ/b5japcIQHo+dTN+MKK/RCPP9OmYWb84ApybgtFaOOXt1dkpRtmvT/DoMyoa
WtGvWYMzDHY4B9f8TWvSpK8BBM9p3Uoci+djWjCcCZHHp+ENS3U07/JNi5qFkw8P
YTsQtbM1N0S1r5kYwrN6pi5r9HDRGb3J+xzEfxwn+nVfJltwtFou+Ds9dVQkN8zP
NKRZlmCF3G7hhN/r4rZ76072Iw9WIgsbH0AblvSgJagal/pIN3uVz1pZnYWsAfef
Hz30xtj+pSzEnv/eqQ2iJgGugBOY4BKiVMNof0SwbX0JOvW7ZH+6RE7lOJMIKtWC
FAOmb2ZH67DDxmWHrnUzQJ7sYpVNdWGT5Bu0WrWXWami8acg7IcdWSbrcWS/fPCF
NUii9DiPYQ8myG77i+DEp1P3EHerZKrdt5ZCjF0ZcgiMH59ItdG0XzHgfbZUJhGj
9kDISAI+V2DLTXwNKWvWwPdmqMSSTvOU4bNQeauntp827Feo/y6dSntoNw7ad9zd
+Msnt0iNB+LbWlt9mcFRuAIjSg/l4eqXaLQ3aeisp1H6cWBzaVYxRq1WXyncL3Qe
xeyP+nVIEG3kDR81/QkUxebcE7+ycXYuYRh/Y2FXiEixR27/wHgaP9uxdiM5KfM9
Yd/BYougdUpD1WxR84xtkurClFm1K5A3HHVrM+ZsHNseCfByicR07Z0kmgEm630y
ZRyCSvGlDMUtJLjAuE363BdskTaoKqxzD1uh/DGH4UidGR8Q5dyE2utdItcjywWS
c8yEB+Fkn0nmGU5lXpg8QukJQxBqn7lrSg11ZynBQ1XcbcTfMscoGRDX+qc0rdsc
KCGUoVVEiKZalc4gPJlXUMO/gk3dZpmZSUpznYNfGKP5U09kcxWb43KiZBbjMhLp
tT0wvISMMMtx/N5BbOeh/7Bkq1xvndDYC+quVaMlBzVE9fnGtQf9BsqfKCH6GvF+
kXZ+XKGg3DduzI5WmrfRvuUQv5JjRH77POv9ki8uqGZLnMGFRmRyXkMVG5FvffPm
+JqndEg0fRP23b9TEWGE1D+hDguBvUuEi4qdzJ0zwX3BOakHVVe2x1ZgvFwUSzoV
ADtAVznxsk16HdJ6G4sp+Azr2pJzoV9d2QPFJsnRGIdfNfHoutFAd5IqoBoprfie
R0nu6CnBXnAST1VKnF4ptwYYDWkcSuGITLYfd807FB4t8asYkTP7oOtEZ3Xtx1w7
fLLWMdS//V5z4RmRquOLIyuwevLkOpOr9trnw5oAewN9eVVxaN5JXhbTH5oloXgL
6bX0EJV2CYdOKizTL0rxlHgotG1dDdcfkK2eTpUw6t+5hDpzd4dIfJeYPO08tTkd
h4bjWHA8QedKCiPjhSKhhFEtxT6lKp8+gFi8oqgVx1k+O7UmvKHTlR1hEzEN/RV9
aaCAuTTcXaMA4DNYrke9rcqnjdIKhMWL5Jog+5wXfrcyqMHQ2HYA5KQ26Yz34cbI
N7lwVvh6omQDQOe609Lb1Y6LuDCNbCsJJ1s4icbzcBUFj427iYnACpheRZM2+Ult
oBxkJsxPBL9INRDGPs8/1EaB6MVNJY5wkiLv+4sj2uLIIusrEAJwnp123NBc+uwO
oAQJMsc321tTCRVMeqlI8uppISZVj3ow+VcZ76AnPxPKkvI2PAKE9VexDf+J+LNK
pj2KAX3xvOirZSdh9DWWYDM8ArfKP18xkbs9JBuR42AY0PYg71W0IGRlWAfMxzvk
DYhC/VKiD6WBV4ybB8Vl3wQ+gjrcR3U6UbsWgvcBBFbMz697g6sLfEnR8ry/WrEj
qndEmbYwW2SpAelNttGkOcV1LlePvUkTdRKobOQICM7nCzmZVrWN6wKwOl7EtskA
im2USoAyOzDgKbuELMkSMMzHfQb5snsq6elfmmmUZ6RIuSpQ3xiCEA5HN0ROUmQU
U5YuZjqjxIWo24bABMh3BxgKSkzQhJ8wizZ4UEZvnRITDwWQGs9Sj4BxIKuAqaH8
5LAEc7u256/ed9KoEYLPvwsU6Ev9FRmVwxT3ABqj/HvWBfzsxfJjwFOB9A2R4n9B
kR0yHb4VLfEjkzkFFG8yGJXY6+Jc3xZwi+TYDwu29wuQV/wCaGOsFP2n3Kr/h72V
5BwxuPbwJVpU/hA20SReuqpnoAms/Ou6EBf38UXHKdE5CzXc1K/kyc6JiHrhg7bO
GKchVrfQuJTJk2lt8NyZaFwFiEZ6bHogP737nmgaqm6BZt01ytM3jOMoeflJFrER
KN+jsMhLYheYzeQzPc+CXxyitEgaau/eNpFgmjMSoaoL44AW6xmypyGF25Ta2WOt
3HT6AVQ31RX/oYFR4v3eC5yDL4J4nnsVbYE+WZw4EpZci26Vt3vXEgnWOIyoOOVz
JCWkYOE7Z5iTE5asssvKzcV7orkFloIdOVc2/Bs1Dm4Bi4cOzqkW/15Xeg1dDJ8F
P+dit7pNl8Vq2pcG3AwyaL2elFg4H+bQcMfxLvwjgo+imMVYv6S8Wlfqds47WPgz
bjpiXB63Run/X4nNqMtmL5rOPbbKrrIrOaivtOwvlaxQYuMH51gErO1EKSq29B1O
1xSAubIlmG0mtI1TOjJy6s0nlGiKiK0+jt5qmOIvJ31U35EOOxJxyiwv1/+zVgcx
Q67PMI63C2vX+NdIPEWqAYB5ffJ3eBuG/zrJOu0jlK6+5sU+OPaF6TXcXO0xVfwq
g3FaS9tIU6sC4NDggMlvV0lNjYPby9al/DHGa+zSjWN7NkzgBzDHVqWZ1Q3Qy85o
SKk6uFt1KckFPlxFxvarEWfVjDX7P7nSR1vVzV0/HNAabTSvV3EzoppYiI7jHVIq
FbcEi+nVH3z0h23LGokAk9hkFxQNKIpYgV2HVvYtqLCePTRq2cjxc5RgeQgnqRjQ
mbFDZKI3KHh8i2mSRZootB/VmoD/bJPtp1BZo/61u9dSbMjBC3sPixWj4o9CJfza
Bl0nib3eTLpcjAPodlYqYpHBi+HHcmC6fZiPf1QkU+aykWXnWFSOo57zLAHkm5HD
OZI3yr3dIIYfdYxmG4uQYix12V5jo48z7R02LSpQYfzfqIQQZbfE7l2ECY2OfbZH
sRCj2yauWic8Hkp3165ugi3d6b677PSMGr+MGhB/pstZOQFBZ2mLNDNJDCaLDhQc
NYJ+/Tyy3Idr4MzWtXhLM2GhNxMV++Ugivc8jx33mS7SQuBmhj2Co7ZF1hg9ifdC
uoLHP2/LXJm6Jnl/JTwDCg5xj3NRfbhm1AMPPuQ1GJlaSNo0ghWXCtecveNmbelt
tFMa0c5Q2MtFWMZTvGCH3OKSoBS92YtJ4WrZkfv1mENLz2Wl8K88yGpARB6yWQZ5
edOAmsRqAO8KHHNuQJcZF4h1p/oLYiNgyVXTmoFPq0vR6g6b1PEXPv2NPv5yhOie
O4M5s4AnRTcXE1WpMU14W9J9NEC2kr0bAyzz1jIwvH/5N6ec27dJM/xCOXSGtxrK
245vJ+5EcUgsGfF+OzXLFPbEkoyyFGZj6ns6CR5HRWNqbcZN8IrzbLxBlO/hHqjs
HQFDPuf2Sut/pGzOfeHVrVCh+uk3X9wdG6go1qy75LnnCEtfiMSQT96WyjSbZvpY
reLqcf0kmD5zFJ7VRd6I2wZTCs+rcdO9331vb0Opxar6WEpAQJRgCYqzvq5TQ/w4
r4KzkP5r9tL0Q3EumAvESTDhNAWgXFJzIzAAN79Db1+DBk8cl8RctW6yomscbzlx
WP4bYlbIxhxlagOXUcVv3qAkPxdYJHHEj0bKwhgYqwD5PzdrWDoD3KHpuBmCfKHo
Z/Bp4hJ6d47LUoQadMpzWE5wfAt5ZprLZ9EyQHUyGuJNaeOTCiSMRmYrlN26yel/
JeAnZw/rVB2yBlHc/TsMBv/h/3TGCY3ygSiBcpDQqqIEZTBHagjyfXC1HqlICIgL
WSuCaaH4vboEiTdLqT7lApF82TDFgljxE/B+Ki1+T5ON/Ug7tdh25cyq2fN40bPt
e+4DrBNCkxR274pRbfs0LEM/xxZKjlRv1ODWE1qQnOiCJMWisIzBnqAeRrCzjsTs
ERRe/zSQxtcVEx8WVtpCTnmLHimFbLKAjyS7In01KclwXlc+OvzQ4NtFIeRQ4ssv
ZBKs6aTovSwBNvqncqfEJpEDdljMoDKu5P49iVIt0uwqoBPChYPw23bf+bNsLkjJ
rDvSmtveYisQrKMYiZYFksVMfTarMVvDo+qm9jvfhEFqn9p9lnjQsqvN2iPNbUB3
A5s76Tve0mLzwAiXuagPAI4QdnVxvQ8zG0SIV7xayjmJpun6CHSMfYXhIPIlD75V
GkxOWJweFs04mShWTavb3WRihj9BUjzB9B/C2bYIWiHQRu+eo90q9jmiJ9xUBw4K
Jcm3JBPJp9759MhEw0K6a99IRdaIFloo0NlPe/WqShkuoLQnAAELsEztJmuMlsDV
DGMR0A/A4N9Ryvtzk/9Cdd2KTT1AYD4JntMfZM/8RKM1uLyB0KI1o8zu3hY5eEgu
v0WwXb8VtYK1P1/K9IMQc8na8FF06lsDKOHaLRKpbJGsi3Z4ovrZN4KBdyQp2uxX
/TNEMM6L9amSwTWWFhHBhGybEA8LXhvog00ryESoQ9Tww7q5gp/oA48NjIK0iSzi
ks3t30rzlxqkeGI2FiftuDm0gGeW6lHFpAjaEN59i07bXmfkLzcQKSpDD/Ux48/h
5XOx9/JhNVEvMF3dXI+K/WID7MKosqgoz3krpBENyawc+MIZNigts2sR16mTEfE0
qMm0pI6hMqQMtwwRKfTKlQN8H4W8pt7MahzovtEdh3Px79lKwSwxiN5WuaG54vS2
pb7WHB83LjwxZIpWbdaeywL9MVqwMnGK5YLK7HV2djvXVsMTOJEHjF3cwo6cIgmk
PaYdsAWSruNQZ4FbklaOSBLz0SEyLthDvXcTZ4RRGe7/LLnxDh4rxyxNSnmVNwTF
mXpWzXaYKB0auGXSFnfyHjM4XONDjyaGjKLbqv2vVdvlEfaeb69w2mO20A4DgrrT
naNMHYQZWdQKjevPp0xDLEEW0R0sXvoYe9HnzuKaH4d7smcXfztVGRGguWxP7wGd
UU6zIzDLR8sQ63b4U8aN2ook5ykRI1rfCeZk+H7vlxdB3f38xqnF15/2x0lp3saB
NM8SyQ21/GiptpCoTAEuyy4QCATBV6OR75YP1nSMBQnDX2M7/pyPCVw9Qqc9e7dd
J4crqyIbVFR502vgr/r23X9pBWZkDb+d3xrm6p/Ht62opvOXs9GzsjfsYHg9aKMj
ZzbeaDRlPfn95gdrEmXqfw59d7M/h8KUfwn5eME77xrb0lxH1aLJAIyz0C3Zc+9d
JSMG/i6Hc4g/C3fCqNZ+wIpOZvriRr17UyycinI47DaU9GZPFZs/cE3QDjYKRRyS
GX2IPQNkJjBqVoyevqwEMbF8GyOI4rXV/Nka0ZxRv/KSgZ2mwheyOglFka0657kY
57aDBPuJHM65Wz6mHmJqsLqjN1N6qD0mbrwGTziH8Q6tIVkBnGpnSG6llKkOjWfj
nfTozGy255h5z7ZQKr7HdOBc0xY7pungrlimMSdfn/ylIlNMdbWrjfSbFHt5ISUB
HgJIQfQcD/1CLkfrrlltmUIjTxdfjW0S4mitjw9ET0V5nJU5ys3+qEKPZgLRdWT2
YSgFPTq+5Pu3+JPkyy5hrJJZQe2r4ztGI2HLy0+LdNsSmkT2ls+FnZYJev0xQrWk
/WCOEzfUl+BWBakGDIOgJVSIILABsBFNg8KqXH1y3wf1UMkUVipkQ1+oLwJ6/1iR
xrs5iETC3lva/GoC2wYtDvS3mYISdWP+3RpdOTfrKzlujiadEkBjDGmN47Q6Mx0R
IhKW/fD5DIH4VAjZXK4NLZOdPIwvxJECoNLbcReI4mI800UIHdVhsyecN1ZYkFs9
Ato8QMfihRhPEEBkzJFzqP4D+E5zetjCpl4v+wnMY9g7vIBbS6bky3nKCiFetrOL
ZQrsuZrVFbCt3WTrnu01O8cNaf+zBF7zlcCIlZapgGdfKvUBFP69rXc42ynzBKgp
aqcCYzBwWE+AJEe0UoYLkA6kwkcPGstet/ZS3vK/zN9vfDOQNiffopwHvEySxr0N
flultFA9s08SdxCIBEN2TdifhzPH4o0yCu2IYQLKRgozcrvOghsyb/IJmq1YIuG3
C3khPMaKjRA+KKOlO505+obSytx7F+3cIADh4zQUkaXF/lNbzcYx36XXXYlv6Qz8
OUACynz8uTqNLXJMdy43376re4aVlHsMUagjSkSTz7aqRfrgiwxM+PHfg4NSI/yi
gL60v9Wb2zUIs1XBgm6uostkNdFjWU5tuBLT3TsLjRSHcNV3wVppePQU/QvJTXOg
3UFIRoMyhHdPaxnEoryxQF48o5C2hR+GME4Lf7qLBM8emEmgaZJiicrIE8qPj9hy
udouh6JwIy85NR5TlBspp9vgEvYihLDXcea1ld96E4zl1lxe3qIVKUozsVudGhzL
2b+ur8+BBuMCM/G/LNyJI30ycWbNDVi0ZIxaaQbCOVunUmpyv9G0buX7jL2RCyt8
fB/JxCxTbIx7cyQP3G6fsH0P86R5uRX/1HvYaEnmO/p+YUVji7ZC8AfzK+QXjzSL
6qdhKRzhlAaVDA5QSRK6Lq3ljMnw0fOTJCC8AixFVh0azCEcXgnKm8PyblbhSiDo
nI9r5ZUSmgd/rE3RlRt1hNVUu+0zBGWk9OePkRDWiZYQTATSU7eykdp1rrk2oVMw
dCehxOFcvuIQRQHuMJ1MGuBx/wqk7rZuonM/fvEQ5U2XMzo/ov/wcBpr/jDwYNoL
guVIUcOOeNGn/g2HESK1uQHsjdo0UnNhc2uhMubUltky5yQgzCDhBRtxLHPS+QQR
VZ+ITtbZrXDsHGxWYsXKApUoDIRByCWiVBU9R+V8Ip4vk3Qx7x/ODsiw1wM2Y2Nc
phXW+Oi9eT54mwvJ1TfIQ6BY+3AG1C9oXmn9/Et0/UIcuDx1rU6ctgPFBE0/Qu9b
wAa4OolotdnvtbmHruJAh7O4ghmitfoY1EZUluiWHS8d3Bnw4wUU4o6FdLGpbEKL
7v9U6BJn1Sm4qyAq/gdUCDDO+N+EArSUK6glO5t1AcZgrGx4agQGFG104PoJEs8C
qqmVJ+CPCX3EAO6sCeM0f8xRU5WCPq1/Ei59K3Tv5TQZ0DoIpLm2bIN5KMdh1BKW
nfEVtOpXNe/RML3ahRQVm4rrlJOzbSObP9ShKdzuoLFxNqZ/M9/BxkQB8s1NzJdf
188k3CQ0XEnrwen4c1gqMIrtVu3L3IsTf6GukjJ6z6UKi0eq32hKfB3GaK0lb9p4
HCojXSMGiFDHfVfRabCrT455SujPGlWkxkQG56JoTqGuXbGdI7Y001aZZ/yVyw1P
7Yaki6scIexSSPTGTUMXrqSTyM/GrgX4W26ao37PJiDqSZ12i6hTe/A8Zr5aYiN7
x9IQSgb3LUDQMBT3XKG72KQxKkwbPe3p3HOXFyD/FHUk7JUBXVxogaNnElHNgeFS
bvoWcQFCW0jAJFjsFn/MX66kcwRPy8nrC8VFADHDxsTIfCO7OSvMRvT7jQNTgC+K
0mSHh11xI3UasfSWoAOA/t4JBjQX3r4d3Qed6g/SJ6dSPw4gSS0dEXSIq8u0fnk7
w649zT8KUeZZ1fBpj/n1Vpsks46VScqTGIhVkrP4TykvEw3wpXRAp30r1PSkrl5W
30YV9QQ+xpyTWxPtGwvlAyKXWEAVknKePPh78gh/DrlMI613wdOb97dc+qOeqEmw
LQldy1ZUpOCiKuaiI70WPr6rgTp6CHRfBZfw2KsFegP9I2Cyf/LNXB39rrKLrDa/
1hc+qzHIdgO08OyDA4j240wTAxqdWh3Whk3DZ5pkWyRsDADwJe2DUr/EEnvsAocn
kJZGte0j7lPm4puCJtrrf7WzlHPqjW7OIKbqrlVAnInFYMH8Vvic+gJcnNfiZ7VL
J4LolKcLxo7a+/ruw1kJPmXP6NqJrhbGHLJh3gGbh0uXzy7TAExNepWCiAmEcmll
xk5dFnRHMgZZ2joDhPygflMHj3eIDs2IYe6q/PwHnLFEaFUPAv/Yr7dEdGldmzZz
V6QMzfYCWufzQBsYUYqSboMCQ/F0al/hUC9p64TETbamlEzGtro+IZZvW7dFr4w8
m3fH1kycLeoEwML6TvKW2F05R/c57JmNOaQ2w3IU9yutqR+Js0OtSfR4mVOmkX/8
f3HQrk1U3i++KtqfsJ3Hn4+doPaxV5ImJKdWx9/onUxNtujFwuCrdkqtL44iS4w/
Cb7/lkaRtZSgROSIK/cIhdl0vMfwvG6JnX6wkK+GkObtpaIDg/u5wRKUPg43tGBA
U/AAQbMMXfpHcKrrCoQa3fkuCQnaeZYGaqSyAH70bJQ2U0FAS6LpgnXM8Muy6+md
188ygEuR2YfbVbxkzydwOS+cGN2qHcexkcCdEtqyQyCigNF1IoC23E+ZtiHDvKzp
pav9EzF8yHKBTY8wRsSckTfmjsvNlV+GXu22yIo9tO8zo2/kpw5rX5M/F0l46+A9
nKsW2Vf2lLjyH+agkkTglqXZTsHwNnKyflmn8sBVvfNjXIv+LaC/jyxxtFYGK7c9
qR37nWRm0pnPda/DeBYFJW4PPzl9Uh/ohck03AJYzZ07YVLKhUAcKQ3rPgUXvj5n
Z2cmre/PbsQRVd8Q+baA5HscM2FROiIbID04DSaMm9yW1f7fHUJgAPNAN764Rw6/
K7ScGkJisD94pyIEH7wMaw5WpZvOC/AFyY3m2I4PPtmrlfR4H9vwwf7eUewUljeI
+xiaCNurpUPoPZI+6toENMLKnkW/y5AJYxazPwgvG7xMBq49KiSKIk8FGiKHi/iV
fstDl8sppXWDnXuFxo/5LJkfjXha0Bps8bCDO0397r8DINKsLngCQD9+sBRmuWBN
A9Q5qb3+BmNkbL1rjXAMAJtM1r8c/CinTm0VJfBSckTqRA+0kFOwxljoPOUsKx7+
XwPhhLM3r+IoazXjnFPs0Qcxrjk6wMDpkcLUoV0hWwvOguS8p6r6acRYdx/FLkO7
3ssuMem14IW9IX+nBSDurvTH/MmmzM02k8NTpT+wuazOsu2PRJEhAO8jzNGtcqCw
ZTI3j3zY0YNzjxoeynJ7qMr9KoVtDT3UtnQq4oRZCQpa4ufTcy8b+ZJ/VfIX4215
orc3E3IRKg/4NPisXrceDJeY6NxVG7KhCBxNSvwhjDNVQDJebqAZzJ1w1YF7Btgd
13cpcArf98YTtLHppaoBFEjTUm/iA6G3NYMYfn+LbRjizfZMkbY9xGN6nxkEklEr
jA1uZWvOF/H2JVmRtUy48PNNEy18ddzs5g0kOjmIGxVHoFpBSzuilFqN7J2APyp6
PKCQ5vehyborLQs+FjBUn3oLbyzPGmz0tBer8pw+nNMZHvd51xBIZHBsgbOUmwq/
kUASoFQt3PMoFFbWcb+mCb/OmzoFUdMc0jQogvAKfe43Mw+NW1qFnlCYa9il+DaX
Ew37n1406aX7y7WUaV0zmAFpEtzABspYsibpapdwSATu4h4um93i3EcpwRndJZTV
oh5c8QncZTesO8W2XTkJyu1SFzh0wNh4yfEXM0W4qmBcpRuhdcbFuv3NdD4jUCSv
9sZIRNkcLGpc4czsPLhndNz+H4XKUStZJ+6vyOnefiTBI+yS4QzZwPaUG0NKY/Xh
jw4zyxeuNnxi3X0Xg50taE+q/dU6sGBWfdr2xKVJxTtvu9xmA0eT+xKYIiiWNYyI
mcQTox3iJ4hitmpQAuEy/KW6jOb5THBhrkBQ3198dOx4hdKcl/xM02CLBuOtMn8o
tqonlmh10DZ/d55yaSJQMuHD+g1Sm2SU8AiEofK3RUWldQ3rEy8P7MoVn76NCRJ+
KgZaSFAxj9YjbkDUjCRt2Gq0sAURLiWocGL1NQffBxorxwDIWUKDs97LT9pSiVgf
IDhrx3nQM5Xi3cyXoLVpb1nLjBy3MplqcWTlJcS8atw2RfXSkAbFyzLhicKcjJBj
cCq5rc56Fog3FQKi+i0I4cqrWYQd5noa5748ETqjgs2J1Si+ZUScJQGzLjshEsZe
NxtFn7/TAtD2MpCWvY1K7ulp85E3WtiGo2UB2k/crrY1C7/U1IVk9uUaGuGfZj3o
Ir7m5nRlG9rnV0EKLJv1GOOvNl1NYA5xvvi7xI9HSdR6zcXcBjlA3RWjdFM+N5Jg
MZz6b2Pks3ygyMYHutKT+W2I5FXaOEuIs8OI98irXMZ5m73z6k8nTVYpOcVrqKfC
bXBbd1qnoTiYN4opkV6TYurTZWRr7+JqS6lH/Ygc5nkuoELbPVgVHGF27+m0ATLl
AFPUlP1BnK4Z5jK6yST3EthdCqlVY59N2i2aPRiHfcGoRKSG21K+3inZt3g580cO
X7GfGWUynMryS4spqyu/+G7stTrGe170H+orv+grY8v0NPgYyJEmtL6zt7TDt8TT
cwKQhvC4R8oZCaGs4/aMPRvXhVACcU8FbvS3zE8z4rqGGaiDkTiz4eJOokFPbXl6
ugdFpps6r4e/8nUkACp5xqMDFicoMNjmWKWhz64kUwL2MwXq6hMiHQeED5ucTHEL
oz6xDUNMpM0sGc36o+MUoUEOTSDF7WKemWfe6L0r87H9v5w5pp5uJT7NcM6mUcxf
wsa9b0V7GbIVNd7Ldgpsx5bF2U1EGLj5ZmtFDldv4VXoaJ7zpwP+aNRc4t+h4Hj5
2LcwhwcRc8ExkwcKfi+EH0SM9CH7ZfdxROHZPyrdld9+ZUJ8hbRlMUWeWMsGZIf/
UkXLZMnbmlFygNkXxG9890NsLE64NeWOD0ahbRNK3pReDph2WAv6GZNiLQ0020CR
yE80On00dfCbI/UtY0VC3Jj4YO9Cc5lmQ2MoAoqMcU+XDeaXC3urauQ0Yd3qHiN2
xLyikYXxwWGdjagWy3wqfoQ6NqkBNe1hDdvue6HRHjRFZyur3aI7lDK7v/fkFXL+
A3qd8QG8xVcn1nJfHSXPc6T6uYSLEaM428D2n1TQwiTuA1HR9ZUNF03rMHXeS9gs
MIGhRnjdQ6jBR7RCysu5bif2dDwdQHVCHLGUuVXzNrRc503EO/+IbC4In8KE3w+v
xuGnWgWiCLty5B/+QSuiFzoWHrkUdBCaooAYGKV95i6PqAMGvseCnvLxQ62KiaeZ
PZvnr0QkBnhQ/pOzLRv06i2D3blXMyMgyz6w7JMBSi3iTuViOtgA79CYJqxAeKnb
Pv1SHJBfnN8pWmjweTSLAyDQMTwrA815IhA/c4D8EzMuSBTRUTkaRCDepnO3ebkJ
DfSGXQzt4w69K0TMy4KEcZC4Y/ZlWFlTpvUgi96zTsPSNvlcOmLcirKEdFHEGgDH
j830AOh4ga3kPpUnHpBdaFHdiprSMCKCRgdayx9mRUII60BH5dtp2SzRwOUykRx2
v5hLFRtYd7yKKGCQk4wi+hqpko09CSsV10EaliFIERvshG09CUeSDSobweMxCQnK
U2xbVw+Xp/D+Hm5tBpCLgQop+a20TVjgtNXXpUYo2BTW7OF5W+cjtW7ynwFTfgVT
J4jyMf6W773QeNO6Cz1xxwyEGCaXbeqss1CFHEcigR/QG0KCVvt1sPLMAd6UeFwB
efFR/j115yL6OlEufLrvBrB1gE+G0q8vvlUgpAdKghkIFAp7an4PsP3qwBHfA3Y5
CVVE1DYRvmfHg2D6I5YgZTkC2WZmYmWeMQ86jqWNUHGgfloWRYml4C7CLXArrlWq
lQbyJ4SlVwA95/UjHd76+dfBkapzSqAyudDOpS3xOazuhVQrY3yW8R6rn2MsrDpb
gJIXzC/P4oKuDp7L6lMHyoIZ/JlAIuR2SuO4qayAu4GqgqLtCnC0xun4XM0Eu1FQ
eY1cZiUDnWSOTQlhdTVx8+AU2kYy29kPq7IOz4B9ZxpWsxszLtP7z4E5+4F/YIrQ
iimIMpnOWZnq287yJ3HEEWbiuBG0MzZ92tPtqCHQMOrZq1fydhyUuUqcCBXetcXc
1l5Z3hiH6yqXhjKTwfiNvX8LGegBRIhltueIjSfP7SQjOqtYf253EcRALjE/L8u/
5aXcnKAiauvUVmDUg+/M2Dn2MvEZCo30eJsbMjNodVLXttPUVDV6BvgY/7halHve
DWklQjUU1qh5A36qeuv8Mtq+bUvwNKj8GkZQzyiFLxoa/hAUCvNf2Z2na/dJaMvP
ogNFcGD1bExAqdBugtkow4WsnlnxSyFt73rNXme6Gzatz+nbg469lqHS2yVls63O
EqHZyp8p7xnprHwJJmcGgsF0SEBZ6qoKVFmRXtFzcmSlt9nusqm46NaFF8unoAO3
UUmHMSa3i7pkpzSmCMcs0V32609gyB53rnG0fu5i1koDafOYqdMZYA4sMv1ntIiI
siyFHeEBKAo2cTpam6F7G5DzhC/p1ntmrrKVvg2EtHXjNASTS6oXZFHhPODeS44h
TH5gto89Rllfw0qwnptBxawsjHOlH9UJgZPeXlAZAbofhNcHnEdJqeqyzjERHA1L
LR8HN6xOg2wFn7VQks9aP7TU99AE5mUfZg+5HAtFSrzBgVK4zYS68sG2S5CS2Yph
ehPZJebIYU11DHpkfRL7W59IGrd+KpmvynabElQP+LmUqFnkrcceHGSkwB5ICJwg
i/VtAoxmCHjukqLpPc52xy3uEpPUzu5QsSrypq1f2R9kMgQi2FwA9nw1j5g7Tp4V
jTfn9m122ZHHJvMieofTj1X8VsgkNykgeQ0BgIC11KFo3jUrHRzjh5pKQSkNRIpn
bRZnMv5dWoNb/lYvxSj/LrQVhdMpqI5k9Ser33yN/i33o5zec60cT3UYfskMN0yy
J/jTpoORJu8gGQWmeths8HaWviLpg9sF5EdH0ltqdfraj33Smp41Ke1BakD4TSHv
3RAAHUjo/NJEVCVJa9QDcp2T2gjh3I1Vd3MbEOH0RBUQhiQ+BTRjkmHg13+GGebc
vM/9QMBDbhUs4CqIzntv8a86i45hQNgyKJL3AXiLzSb2rHeVLIdbi0maVb5Vc0lj
vfrQ1K53UqAJ/Ojc8VvuAYnVPq45OI4DXE5UoL+fm0MTi42yUdcu0uiTu4Wzj2+O
94iQfchjvTzYEeDJiL/8HQAqPI0ibgKVHjaKVZgaw4CQBIL88vB+zx8ZVOB0Mqhe
bpV4+LGyEVNynLQdxQIk2Dd101bw3b2fIEHvSGqr8NePVT33jlWcQfdDy7RcWatB
sDBeKvp+ZPkiFPkysd2hos1BhZqL4Obzha7FllOE/xHugNu67W4vRrwMBbBRWT41
SHm3PhHsJBfzA+EdV/jRYvbYWtlWe4mIF5UTu/9SYriRT3swRu/VP3/K8zuGfI3K
uMr/bKESqQUhD1DD2+98k6USMa//KnWLDm5PCpFViKTL0PSH//orVGguxTV7KFuo
gJ0Tizgg2viEgGw43bvS1Wlm0I8UQWWwf1FPMsqPn9lTUT2DSJBlsNz3f7hDdFV0
rBQSCCmU2i9j6Px+e25QhFmpWCZPKEVAjRKmltOKkf5DKOAdbPSps7gbDytq+snH
7QTysGnGlH3Fdg5ZADtDwtB1XRlSoLTh91FpPbOHMr6E71bj2aVFDpdxRKQO7+FV
2BTx9vgEgbWPxxEzgq1p9ib0jlBRr6y3dJ/619+AVvMMp/C+TSkkW8bRmL/42pV1
DW9K+58urbeCbbRnylue3zWmrPWwJ+RhZS6kHmBGGygYGQSKsXs+wVNy8tgmB6Vx
BWyc/1ti7mKORtthfl7nvrbZ6TT8x0RGCO9ost0ZE5+54obX8bBk47f9M/OUCcek
hMV97uBvT+048lCN+R+S4z0ImM0+fGCGN5kjvO0Q1r/PLHfVU9d5ZpLE9PDS2Ik5
05phtAXzH/O5qK/DYFgdPbofbby02OyBq7NAMpuVpBTPGXj1OriTXpL1ZULNiwK1
ei6L1kAZMuRNHxn3hLdDfLrgLrmPyQAsuoNnd8u0VFEgQ0he9969Ux137OQFxon/
wIp/DlMKf/eMSzTpNnHLuE0v/4rl/E+6AeieoCr2JkvxrezsEcMiLqmQ14XocdJ9
0a9tVWLRN/6YD3TcM3BwI21lQtOHNXthNmqhoSqjkrffdUGwH6+UeNBJ/RPpDgVc
0g7v+FWk6ftyn/ySXnRnbDLDIlx7JIzMY0lhYXqLA3AcZw+EDhUZTqnCxllrBbYh
YJ0KcdXQK9b312iT34R3h6ox+T1Cr/ErQ6Q5ro59p1t/jikEOD0/WIO7I9Wsy5+/
Kr3as36sMNyVNJ3kSnSopgXFlpj4oGQok4Q1a43nK0fS/sFLBJL1eubPt68E9rZx
FeRKEj3QMKObw0pmvvyFX701vcRgkOZYMb9dnvSXjZIRabFte8J/QQMyXmZKjlpi
Y0NJoHS9z2xepcZ7Qgb8Sjx0HzCDF3PlgK3701dDhDv3e2xbTAHXOailOfJxmOdF
yVrt1Yk9lcXNNc5+t3c+3uX4FPxXxkvb5d1BHHpnuWNZ5hcElDOMtw2hsYNiGKFJ
s+joAM0tQU5SvdJ/ycy0+GOM5pTOFqCP7AUDGGaBJYcvndX7kn2BGkisOnosm6DB
SlqSVZqe7TKEYfyxVidCbMji4URb46sB9Z/i/u8+FPrQ8jJCWcINErUFmVKJxL0k
xRyDOfDibnTB360zumtyXfxNI9qyEeW3iovK85OaZ5XDVByx7P4jGNija6mXbDX9
bMJIVY4KmuQ1qBoWypTYulknG3YYvHRBH1lQQWzIUb692LRCWWEeN4xfwZxTx3Fm
uey0MMQmdUXmGwcZrNMH+l7SFgaEvN9DeNX987LYqR8mQMpNglun4yMqOuebuRH7
xdyfMX/8OBrN2hJR3mpkhUZNHOMt7zIQtznQKB/eiMEPScTLhpsFv5XMLFF8cpsU
vN8Ra1+rgO9+Z/3N6kHAlWm//m2vf0gEwhzhCnpkDJF0x2g/eFk4oDbMtvaljhsj
gOCsMKROjKyr/Djfq2gyxBDhYyjEzi+FkhUVQJNQ98mpzdhPUstn7qJ9XBgUKmpd
VwpW34nwnBc/YjVGXRYk7aR3hqScJ77PU6cpLAekfYMCIey3Tg91xcbvDgDSbUf/
VCm3C9Lho8RDl8HOOgUHpbxGVA7kDB8Am3xUwdB3l9UlsisvYzdDDYJSyKjE3NKg
PRBtdNr2wAJT/mv4WWaK/syi+/OMQKQbrlpknmZns3OmhHMrbEr44zc826OwVo79
Jx3AQsjvO+h0ftrx9Ht1jXcKVSfvxVVJT1yLyNhXhBE6RZZrK9Mpy/4kMQZloylB
dKe96b8ww197Sjz3Tf0tDVFIUwqiZFHHah1QTmvhnglXUQ2FYeNlaI0tUA8yZKPJ
ND/LMTGB9MYjY0Fs0Ii/jGRWToZnlsGJI6OcbJE4ihpnH99mE07vbOnKLeyO0lbB
YB0JRZ3e+n8W7uG7awAulmmStjRq9NN0+mgf7aZCSp+nieT8fyJzsGkc1jMgLcii
JHtl8qTbnKe+DhKdOC7uc/Epv1VXd2sit/GSA4Ug5+k4qW0icDkNfiqbHlrX51OP
XyjxJEMmvXndfhl0C4ySmprqubxmSpC37Q7BJ7YnNaXJ1Pj2KIJqlU95cOgaqKCy
vKtoKdbSjssRpbOWleyYveP/AFI6RpXELEThUj2ve2wNHJUPLZSqRPwEVAdOk0r6
FcwAdMvDAjYUUoc74wLWyBHftC0KheOKlvsIEKsKxJLcP1A2GfhiBxRfnPPpwPgG
HPKXss5zhMHd/qTRBEZiuhe0O/a2IqoeoqdxySiW0gNbUkvlzU7zRSuGVrSza3kn
oV9zFLAgevnJoBEX0m+d784YAlyranmhG0rIP3ZujggCDoey7HjflGF+KqQbpuA2
piMH0lArzMh8SMHPJwFMzDTquWglTbrcN2Dt2kuaTsJxdSLEWjQ8KMu6izhJmYUo
dJBDMU2HAsyGfj8Vym8dHhPAakG4K26lu4Dnt9jVjTSMlx5nnQxxIpFRxwjRaumk
zJmju/KrN35X19984UpVpuQ6Dt6E7bPsyR225ZML9pSrBfHDVOgkqquSpK0D5sWy
7Yv2Btw/jmbMFkm1WLb+9+AO+A+WGJQmnAgnzYIdtlqv74t6BVKMFvG7P5hM/JGN
/TEdVry/azVbipwsOtr409ZrJxjea/LEgdoqJcjya4blp112Dq6orlnhgOA6nFjx
HOUdOc/IXqs/JdX1as7QMxKo2nEjoLCm9oKFx4IBD9YydPmlSmD2y8+hP0B8H96J
WLbetwskNvFpISFLeVH9Z7IQLVQJ95arHvO4jS34Ep0SAa4bPefp5ws/ib3akCv6
f6R6Uky5febAagW1vl9lLmyt/zOx0YeP2waY+Eou1gcQWy8t78A40K/+WZMAhSCR
qgdw1IbJabfVNKvRCLRliev87igm5iBh1wRBTDSx5dP3JnyT3BtMplvWwA5Siw1y
bu+a80FtOd/lDu5uD2eUANgkUWg48HLwsJfaZyQLQe7c4O0FDP+r9ikKuqdJm8on
bFD/VRmhcwPQfZXsEzIc4uOM586jFhTmnV3Y+qfOsB39CUCoIiU8K+1LOYJguYDf
TcP0i3syrrxFZy9JUZTgkSMknIffYN8/aDgGB2FvoNl+6gvMXLtxR/WDogzLTC4p
tBUUuksG2N0K/jLz6CDuctIHn3hEUQjZn4C8j34ZV5V5Y7z6Vxo/0XkktTTgPwzA
dDuzS6+1jh7vYZJUEF5YeUOj/eI8Iqnbqam5JTSn7rYBIW+Po8HE6OCi+K15vv9K
NnaBr941AILYcgwByzsJhvJpPnnjosT96a0xaKWbchK+R5iL5zg91YhCjI2CrQ3i
yMwBxYi/Q1HedwttWHSM3HvTLe3gyOorTeRTRbKqP0nEKJnVVV+W9XfxI6QZbFjF
d+JApJZtZpz357ndXaYMtH6GH7BCIWuWi2B2qTozQKR9Q+7BNFPSVDoOyqt+oshp
goesRntHDKWipATkzoN+pLajouMi83PwD78woLKdvbVSs+ZAYhEUKYF5arc1GJyd
cRMIxkpN8gYbOjlDFVE3qrOHmHR4DoSIfr8gq5TvfjPvvnxaKKke4VJLKLtH0poG
TTqJc6A+t76A4yhw+9GGUzWmt4WG2zUN8YANirBx8PVMGBWYvN6pI3yq/QD/6cqP
a/1W8W2Q9bqS0kPn/cHGTEGOWNDXpBMPjieky2FwfuVN9eMMdXFO11j6thAL2gAh
DW1jvbQ9N8c9M4Ij0bV7QxKc3vVuQxOJrzRjOFLKG3tMh/Ysi7aJ9YboPcSq9nqG
sWA3emsGuE1Iqs1P05eErWA8nyWb6JTM5crSv0dH3jxy2vLY5qbXgoGI/JT7ePyO
UWXbP9+TLQTuwIHG705PtKhcOYaxu2D0Z/PEnB8QI88HMJT7zqy7NUEYkMKwZXJq
ymnwiuGYHdlsZmVEoQ07Ptgj+S+q3UED8VK+/H9sUriTieGvAgbncaFX1SBnuuQc
U2nut3dPAXKKwXZ06/9J1/9iVJs0mJoHkD4JnsrOWB55iykoUNtpqqk/QF/YH3vY
A1aYaI7J1pAaMvGYQz48nWpMX5Xh87e9bxSUCMAXv9g06NAvM9oAs9Wn5wvFQk3M
OywltvSycPRozgkFeMeO/5xqImUZmiXM2NP4TEKB5QED5QZBZPANyQ7lp4GOufyD
Vzn0eEI1AuJ/7hGaLdIWDTVk49OVX3q8qPOKZCsbAZtYhC1gYBixNT8OorlvQbW9
enJS+5krhLflDradvxvoVL1QAPV+Fe4SuVqRJhFCvs/4x3oNyMf4hZYgiqGJhO+K
fz6usV4qsGUX0wlEF5//AZR9xUXeXBqqk/ZHEHjsXezT9tmc+fp5RIJTQ2DY4Pfc
OQJKGFV7hprFTa5wnPrqNEhOVbFs/RZ6iudCW4Unv3n3MwaQixwZWIIqlP8XQLes
nwI3vY36H3UyCXcYfiZojwEeQXxIeDaIe5IQzhSfZZb5SgsEnVrNVtGBeXf9fxCZ
TGPyjLzqOYIaJX671r33VCDlIJkYMUl/zM2RrdBZi1Vd5ggEgd1PfPEZ72lcnXeJ
9LmtBP0ivW/3bEMK5hGxINBAujkwDOWGTC9PmemGXc1uY0sphckr/rtwlMsxnXzk
u2TvAVZsZfyxHOuWT9IDTPIPwW6U5PU8iYt80sxrMbQd25FKg7dqlAQe5JII+vDW
viiKIjX5NSIJV3BrLozrxuM1szcbxZt+JPGgoXll+K3rlf6uq/5gBjKabxm64Mbs
Kr1o6xwM9jryRpwRib5MTypOaLRApoydGeU0Zf+OmNTOJwDImqMA8V25BkClMWNo
PkjJ7hnPoIUssv7eICbx47tjTHNOy1Z8QSmLtNiZMBo2ne0x0G9dX7y5ric+sdpM
9fFmnf6MDqT/nHMI8eRvhIdD3Nbh66nw5WyRE9V45y0DppQk1fLd1NPV5Yakqjlp
XD2VdNmwJ4nvFqkOlelsX2VwMuITl0VXMqvIOyFpPAqmFgTP59lU8cYz7ueowdor
DWJMI8i13YVQvGrIbGAT/sCLWNHLRCVVtjChpT9MlwsMCPC2chp8CyDy6Pjlf57D
LQrtUVF6GI8fFqF2jXBQ0BH0bCS7XS6htQ+5ihOe2hwV3CzMuklKAlKVd8b3SAVg
ezaUDVMM52xioXTO91mcdiYvjfZX1anIOc4UFsP2Yd2g3DYREMmivBpR+gtqtb4c
6Qe2wdNJejSs0vmUc6blKuoTEocblxrCrdb6/q+djKMDavHHFBw+6PGvSYSETv7s
cA7ui1rih0iS4t+T4gFlURzq306RWc8B1JzIi4M9SQli+2VB+Fd0jExr+9EySuzM
9ftyuTTGDCcN0IYfPZI7P00ykexIMt/bmC4uG+8tNwV5BSUn8pIZTKFum3B6p1Qk
aeUAxdTQvnHA8sqpa4cL6FM2cwdefY59O6CCPW9vdXJDVVzXs1YU1hifNZw1vz6g
AAcr22gHqaWhwQbE0MveDgybJ3vt8VeNIWw+rGR7kQ8D0UQb8JJNXSgvLlfkXhwC
5ncYlhF95ngRybZkxRuV2KkWZ9VeVXvcisyE3DQtc/q9DDryQsfm2eRD1DGz9lNH
HtjHIKkzPJy9hfHehryviomwTzsmLP1qEarUqg0pKKGNjZoFIML4sLbkrY3fqsrO
SLrO7YQtaDi5wPpAd6qRxgjMhVemKmd/sXznCRueFinIK9i4a8RtFRoV1fujCNwA
7BKLZo2O/okC4n4CzwdHGnAEnMsnxPM5ZnEaTAiEZ5Z9a6ppaOB3BXZysRouF5cz
d3JqcXTCLPhuT8hMePKcQRhqMowaFHPWp62qcE7Jkzs0JWEttcGv8s8Jg96kvmhc
0qNGy56x+/GfxDJ+GypnCoiIkTT1cqJgbDwJ3Zw3UhachhGEMvcqcxf6jMQhnnTv
dVvnUm+GO2PMk/A87G0DVdc/SQip/pG9qqEdcmNGDadolr7xNRkpzI9O+AkeZ0Cr
/1S5dQIQEvyPzKWznG4wzh/l1KFNmZ13MjSPgEjD8YVdBFq6Agq6g0sDoAbAwDre
uDmvDt6IiMW+bDg/zO4MMU30XiiY5co0CGNT6P0EaNubQI7aJOUbSri72dAGvCl6
6GgDAos3fc09KmCF/8mw4Kx6d3DPzJiGlcTerZvU4EkxNONvDvsOtT7Yfpzct0UN
pZhmczmNH8bMUyuwWzbdIp/LSgi/mnLgwBGbeOynylLloJ2AHVlixv7eDejs4xDV
SoG2RN+QOY2/YJUgtox2f3KUFF485czG1eXTWVANTKiM3ghh4e3llyoMpnPRcmGq
hKIjeyj1vHGvixuKdHI1lpPgz7hn+OV8mC3zw3VnT/2eEP0iHtceUZlA7EY/sRwM
PCxR4YaV53RuXr2kVyzu/L938/iBy2GY/wQws9uJgvs1KC8YpZU1H7eemZgHPI5o
zdR5xEEEl9DAVn3Z+RPKqwh8cSdPgQiNr7wbp/95AJObpj7YudHYSo3P8nadaccD
wAGGrJweXjdcPEShXVfrFdCzuCBeZZeiys7SPvrfxVMWhbPJgEV9SgW6738wNVOZ
WRT5nQIUEwicXVoRWbdEzDZZk6aSjxfv2UCanKtjgIlpuE7gMaftA/mjoWMmXncl
bhIfHV/t+SoSQbFWjRCatGwHH+0QKGqo2rhwPovQHolSb/Gen05/9xzSfinTukaE
BSJzOY3l9P5e0bRqH7aXXLaCF7P43RI5Y9XGD/2xdeAK7ZMdBLWpkTd7BcQOjpOG
j4Vr4E4ksDLVVTqeYf8PC7uXC1kslVhsh8rxV2JTTdYXQlz8IuGI8SQy7Zg9ZmRr
OPFu7Kr2WZEGQyyYspEFTacH1CkSd0bLiHXbQPPoPXBXFV55OtNUKrOEqb1j/Ksi
6Nn6Zt0gsnEjSfJ4QgPwEUfImqZoC2c8sF+KoEDlNYbcgGBl/EOgDWcRgEZThsK1
GkM6TotZQ4/IF7ukGCrj6jHePuA8mIPIKXMWdvYIs+q8EwNumXFy0f1TcpjqdV9X
tPsSw6DgNkQxSzdlmqo1xhDLfmJCFjKKasaet+dBwB52t+wvDQmDt5qj/bMVFfBC
RDUt/VyPeTArcickrGNv1SLxrMy1lfNjJUBiVPYQor/700f/u2IV3BO2+b2kLOR4
lJKScLY5t/g7ia1/9Zb6+BXoHIi/yRzpW5ZHtOXHgL32t1BLIoCZ2u60Y1sDgOOr
FKE8IMv03EUvxasP4979OPKcoknDFG98lyEpcHgTpkv5vfrbjzzA+ZxJC1Vzz8Lu
mmMqSGywCjQGa30/io6ZyERzfj59ASCiAwnO4zfcH+/IaTkkqWkwz9rqaQIM5N0+
vKyjPT1CF/gPf3HWOpqzIkkH7q0VYfSSkbB2u1U1qNcZB9Ao37U5vSjh+7jmeT7k
YEfk+UHxGtDqDLThAiTguwMyfF5cQEE7w/SYGIOHf/U1GXKcP9SZdzOnIxPdGCuW
vDVLddyjrKIfCczOZ75+uDSQJyEEnIk09qeN1Zp40Nf1vJlYITAVe1GKKKScSjuK
pILS3VmplyczNOKCtYQCF2Uy/cGQERjDvLkIiV4cdF8uPH5kDvTnhaL2onODqP/e
TpyRH0Kklb0GUaMT0XJbxOQEsNujp8fNZ3ylNnvwexXpgTwXknuwzRf0U//DnQWN
ddPEnfyP6gFm4ECkT6pIq9UNiitE5juofGI4CNCinocKQNJbdDWhPA0i3ZeYeQ+i
HKdM79iBrm+MBdL3muD9AIC3Hi0ZgchqKjVNtN1kojLSypHS9NvC9VQ4Vik/wRfz
pTAZxZmUlOH/AVHpGshipwNuA6ErzsHre2qDG0PkTxYz2KhDnaRd/tg0SIvP2imx
9Anz6ILxGvaYCOPl0lCrVj+KLQ/GfyeDT+wi6Fk0HSlFMahEtDkLjOuv06wwC4a8
nwNEhVhwVo0Q66xayY6CMAABcwTEKt2CIHFnG4d368w9JJ8MIp9dfCb2Qgfq0U3J
3ldb29f95vtnZt7F+JmyW6dpKkrA9ac8K4U1CI7Sq6GkdDpN34MfeqoRbP/vIoOa
AvwuWZSRW2JpdDx1I6boNGJQgqWr6FHZ6OIwgO5Xj+6VqxSu8Tp8asqN4rCLxvVC
2CTGG2yJskUhoVC0LG31aEbKQZ4Ojh8FE79J4++RSJER6AzA/6Y4AKYpsmG1THWh
xViqukx7jSKH2OwHtCbZa8GlZnmahkIg1xUhyeAgTnhG8Tw/YH8UyQwhqoLJ/1xJ
UOt9nSY6lo5CgoS+BEeVKGBmmfeOqYuGuueOVlqh4x9qJtdco+SiHOHODPy7uJjH
a7przz0hGqIZhgbalAou/YudTDCaJwtvisXwRx/LIFxA8gt+gNCmt2yJublizxW0
MaX15jHGyDC3dtBm6/etuZgvH+713ki9VsM3SRQWaFlKViaEGEctTMFC36jtcQEf
Gk7NVkhDmAUxrpy/I8NDXyE1/MbhvtcAzArOGkvqdob2M/gdqr3fUYbLnDdFDncV
K8nIKOdjMeE/RfD1I1vslQrqFx9FPCicFhMNffhCVxTEt4BVGzQKJIarzxk3lNm6
uYn0h0jYiEor0sTKOaC9NPh4KKLDWtjxi1rE9LwJK1q3rD21OwW1RoHH+HaSGRmN
cp0IEk/UpKVYIWBjhw9dNwXnWjW7mbkH3TVc/on3OIsorXsp3D6I7GXmwyXD2rf4
6ecaHMJIPhZ1ctUW+Ej25RzMss1TinGuGwNymula7I1mpQkz63XcfBgaWvmwBSFa
b4naZAx7H+8Cy/N1wiqgi6mlNq3fRBeS5mDlv5zOvFyqIp+OmC1h//3pwhxHQmzS
EwNFXMB2dsbTzCTQIoODoh6wle4HU2Xxx8GF5tbLbJYIjIyu/SNXpS9z9KE78yun
iAuIcu34hCmnkg/34KFtv4ZDKJvhyTUQBVrYnsSl+MpbC8Z3UGK1XLblrRzc3roP
RRHKkmsim8LwPbPmpPVqXZhvTgnxKDcH4NBIy95s8y10Y/vjHL6NveNIEFQmiaal
FZh+j8AzxW6L2fDDjGiAe9iHXwxmCXGR6XmWqw0H6jL8Rm0aKN1p1x68QRLlZK3W
41stO38eGWZ30X8jTr7RyS02fLkPU3Zna9mTn3ekiazrWrs4bAMSC435n11tqW3e
UtsLKyU/P6QLAPsE+BgH/0E+kOd8oyIolzl0F0sGlzMrvvUnd2APoIa8q5uz7NGi
zA/qlGMXI42QYc5BbiSaeGFJ3vaNBgKTeYarUcLE39tpaWUQAFn5scESUVHniFXP
yJ1mROzgZ4r/Qt1BKx58VQPB1qDOC9UBf8uRO0755xJmzX7pWtEvULdx7W4YrHp3
3ie7H3h8kaeCZl5Wg9dD0ACNgYLQCSC2kvMMBV6PKZ3XpzqJMkOKq1MZa1F0FW36
mKFryt5qODEJCEThzq2cb2pAnAIIvTl/uB/8GecYLkJJDR8bDJHyXPjuH4vw1q+G
6XJ9O15a3HF3n2XF82Qf2oJl2j02L13M30bQywNBohHS9HtZs3tA5Hf5/rZXHAtX
Oxaw8/cGMMN8Cxtbo0UbSAsjpCkoWY3nJ2e2Ib2wYbLn/TW3DYJyWRu46blLu8xA
RqVprCjsbsD6JwCmue+FJGYmGsblAcLsABP7MtkfePsvv8bj+Hm1NHYymJ5vlgP+
6AggWGoHFd777E4yHjGahZkKY9yrpot1cWJaMNcpCIJgl0Eh7nF1nySCs7TIMFQC
8phdWh04Az2pmNMGrbm0yfJoVc3P7Ti+ujdw713NgLD+uLJujIzcMYqbgDM98MdS
/aUC/sBDL2Qk2TKVAeBDAdb618hLoAc3NTOiw7sNZRgPk3B2QHUw/zd1YOMNKenw
Uurh96H9/JPpnkhaqdnPAv8jEBWTUnvzXfe9atfrjL+S4ljKPTIR2L+6teXvbF48
ULT7FKvjWXYWCstV49tpNqVNiJFjfAZQPmNCE8p2gd+B8fBX7nA3MHa+c4AEb4kX
SecdYkQ53YU43XKB5pkspaCApGqMSnsUxHgxFFYUyouL4I+fyEhnMI5UezgFzaL6
y4aTVc2WIc96BcN3LmSycwKLbv0qk3xifzkq9unRoLTvFXbIjBS17+PnusQWIps5
MKsTJzVNjadh6xdQoK1gEXu5zoTkk5IlUTHkC1AMW3Thew5+Fj04f/DLukX+/p5Y
ZmE4+0UzThJzd07GbLiqwvVdnfMcdivdyZiRtpHCTSb4VOMozAO3oyNP1KdrHP9d
TICkqc1GN+SqryHuNYL0hsPogKqFK8t++qCo7XmAxE6s6IyQEoQsgfdObASWJwxJ
KJQWQNA2GjllB+GGcLoYPN28IUOHjQoP9ZEZ0stEvsZ2FPwk9qZJJXDbtqZhgWd3
vrPpPlLFg+1MOsjSlAQa5EL2t3AiH8xjzX/AgXra0prTaqLHlJKN9jOoX+sf35vu
aZIBYoziabEWS8eAdEv4Hz6JvGdoNaTNQXI6qpSAsTzHeZ7p6rrb0bCTb4WVTyVg
PCiG30c7+YV3PkUdzyr7wuhp+10b/d93O1WPUHAziZiczsKuY7VNg1+zZuLAlHJY
flSvBgLbb1Hki1sWPGqpN5ND9ViGLZqH3Ie69SmsCzTritW1ddTZOR5VBgQ8kdGO
49R3FvmfoNIpZ0qQT6ws8sW2PjT5qSjCgmhyk0vzA7K7U1fEOQeJ9xNBwEznBQiM
H9aHOVTomb93bvgoSa2Yy8CGCMSHal/uFGFmLL5LbxBawq3cDf4y73J00nZeJLbs
YXpaG5syJICHlz8Bpxk7DqhiGPEiLJpNeFIwiijsXcVG02qHmezhJ/LfX+B/1sYW
MA7tNg1LxzUfDZl6wKZGI1BjnzCmZBSsZMIe497xR1hLvGzklHipD+iWNDI+hYGw
mmXdyyWUXaerBt4yNd1KCHuhvqfvaczBxBX5uT0RL5AVmi168SPWoMWKbJd2nFX3
Z2+VbS0bKQtuknRY1gJ3jhHaOPNwWiBZc/OT0+Z8UIDP7JLuO502jdiKlvq6E4mU
lVmn3F2Nlqfo2JO+f6VS8JBLLOjY3WMMTiLosUgaG/x+dH+98EXHmuLyt/3WFMLX
dzJtLfoajo2iMUlU6RQOtUU/LqXKeWpH6QcM+GVeDroU5Zc/lBQfierp1YXy3xzE
55q+mba4pL0KkpA4kfEBCzdaE1iQtgmwkvxv34Bab+0ZOZpVthxUL9N7kPEmrRj2
KB8/RLfG7uAg8P7kZouIKrCK1phcPo7wrOVufS86po/RrSBz8E95zPXtkyUykENU
eWBjXOqDMCwPaZ4ny2xrbZ6/OzcroL7Ef7g++vZMH9GuJR24ClnOmYkOYh8+uqXc
8bCdl4fFPcqyTVQJoGfSZLYhMFg3qfGsWopLO0r+bHON+B5lxeLrUGfNX8exyBUd
7a6uM7ohpMkQshniwmwQpl1rzJ1KS1SQLuIb6vuzyPzm4au/J1047kuLKnyjUpX8
QYVT56Ik2arHY6MMrIbwisD0XfSui93VAonAGpUV3ncWrWolC96oApy8uTY01VqT
Enl32Leq7IljYOp1fqemDBSDpkSFKKhL6gMMvrMY6vMipfwKGawHwo81LOeLzvuj
tnSP2FfPKZ53RySEKogt+Ui/20UnoMEZkDbrlBdxo7e346uIJNWpNnEN7qRO9HE1
wsvXN+qTr86Cjh3ZmasPtW8BeZmYklvzbXaohnT+UP5iG2pgGbv0CbOTNZQHc0RZ
iTEs1ZuZ+lak9IsTtPEW1mYRkGiGj8L73ea5NdEa42bXcuf7Ftn3RkzH2ldBP56r
P0facAs2c8iv8jHKMyjTK4xl6jQYNZfciWwKXPTDYkt4avOpLMs39hTPoyU/SsOn
KuguFc06GDQzfNnbjFG60LmWIFtz6xj2WL0+7itIfm2OHmovDPA8ezn54FryzUPR
U0GdKlpaFg+nnrz1SBNWsswmupAp+YQ5UtV1OaijqBUFOETGgyLAg/AAQNkVQIGz
ONBHB+tmCDnr2vCL6jn6ZFzK8/ClrUismKhVmPPstSn9VAhvFJrzYJmY7qJid5m3
cTkbyhoH6v7D7IlYnRXqxvKZaDg1yBybW6XluKfNHvydhKw111ChI5zWLqZ/UhXL
ceEW773/E0QzjvHXY1BqtchjOvVQY+u0o2S82nl+Ep/ag+qM9nobDxArRKoOhvfv
dSkqiGSxPAqmu3Y8/o0XiJZmck7cwA+3r9mQXZxJTZLTDfdJzm3XRsYRMvFLK+jF
dtY9ou0qR6YCpGbHpZSg1zekYID7uOZ3YnVMFlnMsr+gD7k5pf2w3SqsrJtxvuYS
9XDmQkeCvVQpb5t6121OGn5i6oXSXsQYOaJn+kd4oSOPmCMfTkXdnV5C/Tqaa1zk
mniRyYXbHt9dCX957A05JE2VudoHBQhIi11RpOEEz7ErZTPdCsRRtjRsOpjknLqY
pqZSuwj/LglG0sFJkU9HKT0/3vBeg303Md4O+s/sPw85C4c7kDpYn8ZyZoJ+HmqX
0MslSNl4NQpdrBo886e18MdAZp0iMPrrgzRALRHMCbneILhSfrF6yK8t2dJstUZJ
SAtG4nUZlQpFqYwnZ7CQZU8AxXt4QcpEMus5K2K8T3Ij4Ptrws7wpfkl5EIq7E/o
CFa2wJY9nuadjiFA22wuBWsi/JFjTEM2YvzQC9xXp6W2aDW2/d01DqFoOtiChHh4
pcvZbcmfVKzfQ0Ier/X1MoR1VRoptsseRgqhoysdeEkBRPNNCiif/sq8Z+z+fBB7
mVRzCSAKs7gJli2Hi/bD1+OBa4rJUdVmsKkAAUXbaH/qQ+H4yjvOQKNColbkXqni
/SKQOb6/air+dRszM9N5ct8GytepojNRKRotbUV6YMu9xX7SbOBdMtd2eDwfCqEG
Oc//jeOFmraceKxlMBe3mdG5RcdvmgFKmJMqfLcv5UiTYqJs8zvnfS2HYsc9uK5a
XxChZGEBhjwCSd1EIO9FTN3OLypcD1XFWWS4UKLdZZ4zbiTS+YultaaZPqAjc9yZ
ovOBm0tdwFwRHEk1kcuvh3HiNyLylgnhrxVAavlc/6BKsEjscBVoa7C4ksnReuBy
xiWyIxt++2bl+tShFwr2zRzdDNrrR1HFZMnVVhEhkQLIWqhTUWFjsq4mcxqaa7T1
IEEBfbPqMffDFJ1gVlzzJRjuQhMnZePaV7JDtpAYGwJG+vTFDM+0h+QlgajO3S4U
SpbkC/acmlH7MSDZ7DpUaqf8bbNV4mJeZPNALc0yNtQxvzqvL7Q6tT92BQSjS6e7
6P8OC7fhgAV1zoJ+L3m7erBn4uxpKZk9bA3SDsl6qV3+NvX/esQqZ7xN7KzDcnGM
bTQ4rq6TMFzNQEsxUPSO0IbF4zyh4CCVXVAwo2dv86/H+UGee/T0gS24W5E0Vl3I
VXbK+7p1NHEj6OD6mQ+pjG0tbxDNgO4R+7R5+2qtaaWBWCWh1Es6a+1rCpITmLP3
deDOVQDIN+2YjrRqT7UV4JjayPdwIzXd26DSFTUXrMQZbCPGF36/UcHhNtRNX3Zo
PKqiELe6toPC5owrdDe/PG31LU1GElRvpG/bxW9JnAUjVki1SGkEC5cG66naarzv
hvo3fI9c4MO6k56CAz+TELwgcmFxxn11HUI4CAwQFwGKmPyGNUZWqOZgdXdeBNk0
E1LR8m+4Y5FjNyKz1Xkl4R4FNjVg2xKBJPzGjypSGfmx7hUSWMbt2TuG9FVhzUot
VEsLw5D+ehp8tMG+TvELAqU1DSO9sBs5+cQwv9WguQ9F24pM+sIRMwhal3WUZFtA
KyX3C7ON4s3GTD03Gq/JfaOjfdf/GNuMnNaAYRQMxO4H/wsn2tHuEukoPYjHZRbF
c0Gp6r3O3jNIqbWPLujL2qOc2XMGeI/3BEB0rQxS3/P6B5wCVyk94karCNyd9ybS
QfWrLOzt6GRt7mL7XuluulUGTL/snyVq8SouPJTRT4Y2GyD9VkcyJnDNWsLyVttJ
4f0ClX+EqgrHN8GlYADVAluA7CaWlS2JGy35nzekUO7ijB0lcQ6SJKbjrh7u69Ux
9tWSrA1yHqUppPYrOyHLi2Qkc+8zvSmQIpSwrM5GBYB7JcgeApspiIMnCf/JsXsr
0/EjxjCWc0hIWizAZRH55OYiyIoUC6Wf8VKVDX38WlolWwEMzXEPBZ1355bOjyTr
W9hS83Wno+BhwqzCPEpQpIs4pl8U2K3NAsrvcrO5eBJm0CToiaD/aUs3K2uBW/Z9
tDYCXQCniXAWzPtt3HZU48YQvOfqz13a3dvYY26B2I3DADs63DUQjEMD8O6JbDMr
vf+Ypb1w6qOMcfQmjz3Yr1FrFrMdtEJpLmqEbgbif5Ialugajz5bIcZSakFr/U72
qML9hF5OUOPaVeYQahCwYkhHtpoC3nHkIQNtLBpaODQQlr3M11ivYaH6LZSOKWJh
MZvMKZiE/CMDCfvCFJyw2/UY6exyImnQF3NVnW0uzAQWIP9dIPd4wj6lQBWV4rYL
nrJqaaU57Jg4dRDd4HchM5CzAOW82cbIf2Thtw4cMY1t2Wzctd87dgj0dwQ9LQPv
ztwFif5SuoLgi25OZrNe70bHxWpFmxFSAMu4s/CujukbSVkEjxp52nEMUD4Rukvq
YcnzX3YwDxfn1ki8MpCqAzs3QE8Qykm9j7iVWEg6slrS20eWPixw1fFNwubq71lT
W6sXc1VciDZ748fFQFeiqrbPE07Da7DLlw5WXblhb8L8x1XvB7rtjUrDZpoITaoT
m6hJTyt6MNEsjcKBzX1tKQKTI3uScd1pTaSiWRl7vJVtqdMUYNd/WJCljJ/ESjmd
oIGGHROJqB3o2M6okzPxTaAuTvd/Y2FadLiYmac2QKsl4OzrYEiqJzUDdIL/287i
S1ulC+F3bCLCqkeFXFiYEXnc6Rx9C4NRBH8secQpgnaSH8B7PVsEDcV9vl2wkwHs
4/348zj4vdf07o0wTedyi8xQxCky/0ax3/ZeIPoJJt3jsBxlQjxYruNRmE0AEKz/
YioIfcN/8i99tmcR6Nwf8zJ713SitlC46G9X0D4bpfjSTbw1oUFxsNTS67Y/cqJi
SqwypbsFB+UkgA2KrK90JMyoxhcCrVUcg74Dnnvi7scqfxWEm1/1Xnt62Bups+z1
H9n9kZt3klNbI0Z7vBOL5du9pGRq+RfVskOZOejrd9mhHAhkmnJbq7i5KzCFQ7wr
Xblcp5aMH2RhAxRMIDCwhWiiYZqW+j0TFGPyDFhp0ZuFoHlYjp8CJ+SBppc5mp8V
PVrpCfrcbtK9gfbCVS4l25A2Bh5pxXpINmmcBEGGWFW+vfjJpv9arbAKNBvjoHRS
pT/yaRvCs3u7HAUklhMUXURg4FvcxjK5mJr/2GiBRB6r3QowJ6vAkPL6B/9PuPjZ
xNUvpjy23iPABgxfarzEEDxUTdr6f7CmJB9hDkHEVIbieilJbbvm+Y4oRKZsP61F
5SDIT94qLD2kIOotsbNM331aj5hOFVgZfuqS0n8B4XkdpZSswz4Q0czauJFd68mF
jcGvcNTXu43UyheDbSG8bMLeq+5cDUXqe3qHPtLAdATe3wHXk9cuBdSR3vqtcgl/
uEMOsIDTqZ/N0RJ5jUAZqveQfD29h9dlJcDkrbzZBoL52lsTgRuDr0JazJrsu/cR
C+7Yb0IhSCBh2fXvP7d/S86XqJoIA1nEXc3KU69PEfnGblrKOxmEC8ku1t+65KJy
PiRxZP4TgJwxQSzmnwaxkdOv940epvxqlE7Lr38+08VCKBzWVfb7gFpJQVa2pGi0
eLRC5wI2vNfHN02eLcCmw7ZaFwnOTf2UyOGKnvGPXFQzFv7g442H4nYk7BHPS3gR
Go4y38JySM8FZVGeTS+W3dGHQDeQ8lFn3bLQOXip7cwfg7WnxBc1Zv10mjP9PZaT
rvjJBZhZ+6m52x+DC73T8czUjq7XAYvsuMHgp7k5lGLDPG+8rSKZawq97Z60CJ6R
tNZ1GXqNPieMrUC1L4WqkWyy7qhMEaGv4TFcdw+fgRlN7MqPIXpD5xgh5zUTXQhe
V4iiKdMaGpKqAtUxeXJwRdGAEB/kruDOAZuZlSObz2IOfw54cByn88DovpKMJT8N
y0FYr6yB94TZ2c5hL8E+T2YdEh1U1exxgBRFdCt5IUGJAw11et/96wMssRqwWMXk
rNeCpMhGVO6FPC6oiXOO53z1Z5m4zLmXtHWMvGkfaC/mUnBtdfi6nP670qwAb0y8
DSm3TUaqENBjoXz2xRlXrq1kdZFPUl8RNEArVYesPcLOHcPZ0fNOAEvei0/8OyJm
wKsgU3b6sbjgxswefMQQiV2cabdZY2ui9DpaBGbb6zD49kenPY6sIedheLqT8cAz
pobFY+Q1diREFGWnUF6N8eiqrNE0DJECleWL9BTzg0G5Cbuf10vfx9DTfVmMem5F
U5nwsmB2ZCcUPvgkhB2yVwfnFmyxjMMmpFqhmocdoiFkGP4v5iNLwMdafnJyF0XU
s0h+ljGRVbvUOjocFAwNO34Ec9oCq6hauhH3BzzoNjf88USRAAcigbXX47AjKBTp
cC4EXSxOlc5SmhyAM0muAFar6dFhAcUqOOu7g1W4dJ28odT0nDzzPkYDLD5408c8
ZDU5mCUtwTmEEg2rZ1jf9ru7eKSS748lllbDzxhzFNxmBE2ZC8iOfgzSg0LR/l+4
RkyMA870tae1Iaf0qBhhFxPwt86/sydZzm+sdQRQ+GRzef12igZTM3pKJ0NqanBk
gevFZClICKM8ZGm+H0MJYAN1NJB36q7DdUXLdyro8xvNXcSigATE8I7xvDWn09iS
QJE9US8mkce9h2dAr/6ddx77+jP6VT6iGJiPDI9iky7x2ao94H2pSVORfvWQkArB
sOudngD4YHHfV6l9Gn4CK/xisYAkp3ju3ENJjz/03TxgrT9ufxUHoD4kYwnWGslP
9ZWYXRT5XMVrTqfqm/5PnmLSB8jDJpoPhR4ZL6drIs8hGI/1tWxZXpe0Xt5Wg9VM
biK9f+uTY4fIH/R6rqvpAMLb3pX3rt/YqirSkTurTsKBEsO/3Y8PPds04mxnAw0f
g+EknLndRkPrJY0hniPJdaDKXxvIuJXRG9uLUQpdecSGkG0gJTNCwu1DZtuiO29w
MnCPyqfnhH9OpIy3cGHLa+vPd1Zb50FW4hnqyQva8LVsiSID1aXup4po7B4K45SY
RnC3dJiZQfMhPvqAvlbKqgMZZqsXPY1OBqSG5/BWPoM9bec/jU0LYQT3U4yKokBq
XaeXsfGHswFOKnw+OdWSfl4tKu9tlSCDhTzBMHTxYaDau7DKdzqRqkmzJ3nCWS5Y
STl4S319TAp/MfXhEaXGc+7hC1NoIKV1u6EOBcdzfWd0rtESoDO1m8XzpRkyu4J4
zOf+9nExpLziOQtylS59zA4wKwYZlBKQ3u7O3UCXi5vWwxq5CInlVs3hb0KJPrZF
EbgaRidZhxS63cKtQr6tX6x3M1Y9BnXCMdaaHY8/VhKODxHtVTlmBHXqOEAmFgxt
VfIMkkMSaUoc78kDTGfOjtqb+KXCwVeRwyCo4zQE5hBa3E5gwpz5RpoD6SdPlQP/
zd4RwUnzIDu0ZWKWvgN3Y/sHkVS/CyHWjXCecYLbg+gZQjEMxHxhG0vgDeWxNCJr
u3Blco7roHRV3SoJCq1sBjG2UxXZ/T1DlN5rkMddPhhH9VltKlLn6c+SusYMsP9x
pQ6OTPdZqmcTH3keJD9JS7MwomjpTeN+mJXU7jdx2400utXODD1YLLl3+8JTgM8L
bcCwAmBpr82JuPUED8/cELUVbyPmR8gp21kZ6xqJ7Hv0GzIEddI8lRDMihpKwc2z
sytSmNgJCkuLeVqtE1zMvmkFoMMiONBPj7SczyZOfo/+HteGYL3UYtYNG3t7o9Ii
UvEBVNNxgp1QZUxEgo15oldNEmBA6FJhhVY0EN2Rl9mmwMuiEKDfV4WJuO3fSKfs
Y6lIkORYg1slLtYu3cEzhCm0DV75dlpPlsACv2plHKDaQFAPSAxNwCbF9wSVCpyR
4AKUpcZY27oRAgXvz+fTxDNJGSHdqpyO5zOzj76d3C8KlbtOwPqg+ywqI/17oDD9
QeVw18aaaOEKiNj8YhxkZYDxEi8YrWY+zHQ+FiAEB/WPQmEBEhiq/aEsh+47AFZf
L7qFRpJacvzvf2Yb97Z6WMTUDmjMayxzdarobQvFC8rAii2Q27GeGyc9gd9asTYr
5X9C1gHcundk0iN+YUan45oMh+sNQc9byS56XPBhNIzECTS36j+3jH86QSKNAie0
eShe+bEOJqoGvRrwiFzuJZGnFyKN8KHmHx7KtVV8lp3h0eB/oxSmabVEPMDusDeQ
zkKUVEkayHgJ79qWjYQrG0qvlavgStilmlXs+yjDGvsRoH4TEXSs6kjmyL45j8Dc
KEOQ88CBD2CAa1s8WUcdwneI0SESPoNFByctbXDp4Y232gIan9S4XvPfmmqQvYVN
sfJyOmsVzSIeFnZKjumOiPLoxH6gW7lGZYxGEeATmTCQqCCJ98Zo2qeIT7ARoFo6
+0tD09VgjK6GAEPXjxIZOSdoSCIPDpKaWDiXmt7326cxqAhztls8qhtmgLc9e7dL
Tn3x1I7e7kcaBUeVRg9J0YDwVMsnNzRYPYjdoBRK6ZOnpoluuu2OD9OS5j/VEcXh
wkYb6bABl93NUEfFt75WOONq1sTpYYCz7+t79EfoPN5xfEhQvFiLggGT00NhUnpT
AcpbYbYeN+YgA/3A1Y7DXvMplMv9DFt1JNVZo5Linl0CQ7oKnDo34WAJ4o7CASZA
Za3k5dtfWDRie+pudlncZ21vpIMsSp6ayrlAwj73PPo++x53Hkofin3l02zFmc2Q
191KpU9s7qVFrhF6YSMXTJYMGqV7ICUW/HacbHk1BlwJx125bmsOfOkcw8Ov0m9H
cI9DvV82iKwzcrF+k5Glh1WG3nd2ZdjlaJcT77vAGeqzha8S/JZSYjTn4zk5GkbJ
og0PgyQH2aGxoKooB9sjc/PtVGmT91djO22FVziZnf822wzIY6DOCNDDFJTie2vr
qGSLcSKgia/g5BI5is+iNdVaSoqTXNGtpKPhYmem2gW6wr9YcvMxPkDcYDeowj4/
+cxm+PcJ/0OSM3kbEZDnL8/293jd6fsM5l9L0DEpT/1wLX2Z0jOu0a9lQ3A1rBvQ
P8k3Bo/Mcj+KGLEuRA8R39Ri7ZKHFx5Orv2Emu+IScj5CjrOTlUG6caz5cpt8qX2
shmyaYccUvFe3hlkuR8QcRTKogQ2QK2n/LIIr5isPq/SXVmArFVyB7jMhYkwwkUr
g3HIwJArLR+QG6+dvZGygi8V4w8Dfq0sPiJ+XKoUt53G4Z2hzbp4MYNCc8JnNi16
9QHOWeP048iLKdqHQNLCFWDR9yn5wfqdBzxin+JOg4vQXpwmEb70ISopFtx+J3m6
RMOk0c0X3Y+XgdnhE3F4YJfha6bnyJFZFv2H5BnJCU1hGNHWCacIQLZirCHxyR+B
g3cEDTTKwp7Yp8SPTEvmopxiUgxeuwQsvfZWBLQ/oqvUXTwmv3ofB9rooCT+cdDY
ylnTRpa0oEaafJK+1XE+5ma59ijkIiTg9wi91Lt44UOdKc696jsY9r+OiT+uoj0C
H8syKFgMY9ZCj+whyCYjJOh2ApY12vWqiSQmDlMJ1aJZm6GGWmE0fvNOLVAfvf8O
h1Em4BL9a+Dsbp5NEmZOK+l9e7WLO/zLpiGan8Jt9crokTxYcgjgUzoMh3UHlKXZ
jYwchqj/cTR/WsNrT1Wu/xyXoz/YJavMlv57sW0Auun3sryDhmui+xsCg5ppljxR
QLiXHM94v7dP5qA0cJS+N+ekeYTNsU7jwfAqP3JqQdBrGgqEtn8YoVYOHyNw/D8y
1+gxViDuNOchVR6+wUXOQhaTVe2aN20MmiubEN9HPeqGU5NpZEBLW39jt0Fw8IiN
wWJVyNpBZwj0+FXvlJTp5kiQt5xQb01m8H8sXMUaGdFTFebcP3EuIESQUSVWrT11
GUmhtqihEY9daipFiEbG+bbg3kztHEdVkvPhVv/whFSUeQ3U53b+GHxR9X8tmN+P
om2wC1wjTVvnSYvdR/LVrkAcYr32zSUY/dDZOAKHQ6cS50ifS/kFBg6R9QjcTKfe
bZwzMesSvi1Mq/RC9ldqFiOUHRvK6wfvwpCIP8gf5kYKa9tRMYtnkETpZVITac85
y0a0ch0335iRXCXe4WhVTNXsobsroIRHzDF4P+HxJEM1c2evAxi7dW7QqFmZRv03
phevEpSdojL3cjeVAy/way9k4TLYILtydCHfAXzoW6dTkIZ4lSdxkb/ZMfoZUbm/
QycQGXj5YWj3usbsPNBZGbcaJCElPOcyGKoXlwfcmbWR0PmGDwEmDprMcyapMQBE
izq5XlOtzZeriMJiQmVCAocFnhs3ny8A9I7YuA/BuWwnirB/pO6/7mjWRNN9zo/4
Nnjc6qT+zlh2p4sxPLEm3My/o5E2gdlNUkND/0eA7cfcGbJdX/gw7vgT41ZeEJxB
4egS82EqGFbXVY+xQlYapGnKfol3vjZCD71Fd1ZedahcQeBNl6/vfOUUtF8z82cq
oGga9CFdfJha25vK//8tjtxhWwJ5b8lx8JE6XJYdJxa20hgqucW26j5ZyWOaKhbz
7bCT2ePTUv8JjJV79xQzqd2Kr6eQXnsPhQPYd5r1NiXz7oF+90/9gcqieNoYaHqZ
++CucvNFROsrV7fKb6siTWPA3CqIH71ltn/b2LWsOduFuLjAnWDts3zY6WBv3g/l
A6CPta8vmry0LAS0K8sPeW3xr54GWmmbLYFQnaWfz1nFOUqzIO11Ycm4yABHQ3L4
22eFk+QMT1cEq+dlzsA1a4s8BimQheEtB+dcks95s119ytMwKLz6xGfhYCihs9+o
Sg4G+30FPe0IHMtYm5fBvOaQGD73ot30PIc4DOr0YGZHSBT+iLZYqUmllsBgEvag
74OuUVQqIZI42PbbIhKUuk2bGqMayzbsBaH/6n18VH4d9rq8dZVcWv/pBLJP0oR/
b0IxTsR5G04CrHSE4sSXGzS9vuiePbajHj4HUGAq3U+ilhDhOB8ljbFFyX6Xx73B
jWDtkD12vnb8Nh1rBzuuaV59JAe+oDBFmfLmHCL2w7FuZ74q6d/5obpqGqk7fTHi
MWkt4FtZsUCurRBWeeAAtVKt0FN8SZZEpMbtGPNTbRcHMZbzKICWY3wrQ4qKB5vi
rxjtmRxQ1NSC3WZc5hleQwhsB7t2gPGLBOdTpq56KiXZ8H7K0lheVYtRsrVQum7h
BfHeHK8WDLE7ENab01G+sYmeXfxFKyiNc92dpZ+e3dP20RXDC1KkhQ3JfzHgFDZk
FfZbaqeLCLnCRT8Zbqw1gHStyrx+N7r6mCEtnf0bNvJtRfQmpAnelCSj1M9IxO8F
0EW8H6gP9XOXH5agOfAzEWJYQMqAZJs4+O4p+OHpKyP5BP5+X78h/Nq9ER1PazvB
MZl0092M5zA2gFWKf4pg7Yns9LDhv30sfOtf4OEmwa1NDpYj+X8PWmHx3viQLtR/
c8V7C97xFH1h9+8dUukho5OyCg2UitQSgEix/8VrgtOybeS+BHJFzbpvegjavTPF
7XWhk4vbKuPhGzkKWtvY7i405jSFeGnOP15C0AdD4KImoVmyfYUUhzzyl4GlX2UN
AB+cLkbvE07L6K2Kg46udE+qfaMf+Pv6ozOBg72sXh8VwKP+Yi/VlEYPk6kJUY5T
jCn9eD5/NXwKu3sBjR9fMKuj37v+MvhNHoAJrEbjg6Zw2DYHJgO7huzWsKojxX+B
6VDlCi6DCzy9IAJIqmm2LYhq5eWSvQC1M/WCQxq1PDWHJAVgnPlXUq0b+B7A3mdp
TmBIOVPYmX8f8tErkWo+7aby56xgbEhMBxwglW9frs4tGXasn9bVn4quNO2cx2Ud
MjmVV1smoTi/PMIo2XuCIRFx+Z1VHut4he1BnN+JFaOfX7uvdRxFdPbCe+zByqqb
7WiREkaFPxYPmW4e0NMQNTkRdKax+wS5L8IFjqGsbqmaW3EHU0Xl2/h4GT6rHWsL
gSdQbg6JcJ/f48A9v6c+p6sbxykpEsITLj92qOm4EUfH1ew7c2WtgjyeIBh7B9SB
dREgeFJPpK+4AJJbp4UNjqqYyhCEpxWsZIjmleIFMncUgKoGyl9/pbQAygab1Z4b
kWvhJ7VU6c7YwEDREcQiZ6wxTQn0Km5JAucPfFxDNVKi9kpa3hU2QSJjKgvaTfjD
Xei0N6l2RjU5Acoxg5o9EwVDaVh2dKmMKvn6kfBI0zLrAv+YwOJeyP3FwIdg+cgI
8+3qMqRcq/ous2uYFg3wvcNfQzHHoQ6MeZMjpj2r6fk8HmOFk3f4tDRZzh/nPQ5p
T9plmxMc8IhXCKnRPD2RwWeqma7sClZkAwBSXUNWDLkx3ErroldWXcBuMYtanIXm
6ME/R4CzwLp52LCG7WMpGcNRAf6CJ/8TWTjTstnjkAOKVxzLEmqhzkuQ6lyZNL5q
9JABZIM8EVcTGmyVrW+Rjcv4NomdUdB3CQ7VygOIlFsdgZk5BzMSlsOXI8NUI6oE
+eiachBF3h4LNo99QHJGxhj/1ksW5so5tandqiTaVz3tikuEwAvAEQE+/LSxidZD
Yy3/Z2PiGlu1K1QjUIGCnWwh7ETG2WUMQZyEjoHlqStdenR2cW1/xvKHBMfbMXtM
qjmvklYNMjr/mYEP+6FO802Rv0hWebXbIbiX90JntOIVELgzFMFXr4p98j9yd3+f
BKRmGFAN/wLUhEQI2QrUK0axqZjJ/SOk4wrrA0UZmLSeQUhzUIkV7u/81RSD5f1w
tx3S3prh4tB9KNFh5TPIXe+Mdu0f6S+dfMShgndlyX3ZNoJ4RrI4ypCHEP2yIPC4
JUWm0/HwELA6LtpD9sWjsSMsxz18wX5WBtXA6iLN7KSq3byVf+ctA6eTlAWlMZ0h
BDFdc0ueLAuo8Tviw4fjfsEF3s/rzosxBUED6ryY3ERHTLzm+H6VcsaJJ7TxSazf
PpONI5MhwPS6lgdel2Dh3Vp2jCxUdmAfcBzC4/NytV9HI7fYEsIA5APWlz/tgIcf
rnU3b5MKMDp5Ww2IIHSiCrJWkt7ZjwQotw4NuFOmBOXAKvpxkJgyEv9TQh7t4BQg
eRzGRnSie0pC7ulPN42fgT4tEK6aLEUTWcIcgmzjnovLFagrHNwIrGVaFELT/EQ+
itqzxOma17OvYwzBQXl1VRZHv2z1X7zP9iJeQ16ZpumSYemfg6Ggn8kLJ1UC2BX8
kA6320KaRYNeua4VHPe0mga0Y7Oh/0tKYNR2wO6RRtwzHn1JcnpyBYGdZ/BvkLnf
T5zxDot/OSdzvN3Xn4K9sHFiEUdLWSNR6okirxNt3mRJtUiiyGCDd3QyfwCociWn
ocMCdfCGFTxxDhZiWwCf7jBEYbdKqH7QxypYI5mlMlP661tJxdD7b5ezEBPq3fHD
Or4yyfubx0KkMg7/jS5EUPZbe16kAYB3P5tBnrriYTFg74AU/1MiU+zpbja8f4nc
19ivP23d4tNqyhj9/S1pEuso8j8nRl1r7R+3JPebf7u+rCNsJwkxjZhaKRvHH7OE
JWlz6PWHOwSWP6LaipUhtcrp/HUfQnvS0Gzk/mcqO10YmmjuzF+Pntvh4cREKCit
FsoYbCOc2ZqdNrINxBdZ/GltLs6mN/Rag9VRzHGfDQQct0vBWTRTMtWzQl+fMWPq
DChWRoX7sDlAz4s5Sd1ZXkEdvaai89IDXGXPpjRNgejkDtcn/jG7cPPjpc7tCeZU
A7tqpKREu97nCuSOYDP/rlR0VTYE4CT0BaoTMQeeQnf7LyUv1yZdR+JfTPJFXmXh
8zi/rTBwuZFdV13IED8mvbmBofAVXK4peTXawUN+YyUmFdjsvyEG+/kXYoBszMxG
gzxOmdhNP2lfCFuUs8oQ4f5xURNEQIpcix40dfoCzFVkPil+RoZNVQKjlWDRTo3b
iox2gXjVoUAxLrfQoHFe47sBdbZweVfgmsJoGZDIfJsgJmEGBxELOswDtxrYg5r6
t8rgzAS5LnrgcPtbOwX1w2kOMuGJ3UpiKDD0KAupeMVw2BxB0h45cbUQVPWESzpt
YIbYVksDnkRLF8mDamgN6bon+h92Eb8NQVJRZ9Mcj5y692Qquv6eXkKrRjMw4N/8
SZGpqwN/5DWstyKXE9QtaF6Ytug0d9Vqkrzpd/Ad71gW8NzNk4YYXXHed3Hpb7jR
33/uMivcmY9GPNw8SD073P2pQfoV2GwvjILjAerrz4bkOsQBJPEO4nOvdBSNRtrP
zauCEqG8wuCTbvH0XKD5fJfT6HOITVWPE7inYwN5u7WjfgFZcRNJv81YfXBlcwIB
nGjRs3EaFjXXE6kiAzcZ1P7il4stXMHe/zYhilXY6QYaEgOIJxHpOkMJ1QcKKOuV
1omc5lcK6e8cFDI8cr3uReDN4AnLbzcFh250QH3RFkh3AxplqYgjk58bag56GcZB
J+DitWMhMpCGm2oGcSMau5ctZXqOsvA9yrh/lWBS4b0WDa22OoNYevrNjG9e18fL
ooFypWeLA+UJbJ69wHH5SZM70725BuesIsRWAajcrDYeLU5O1ee+PZRVkwERahQT
Sp2Qz51ybGFvnXRvvjBV0Rs5G0mAkdqyODfvIQFKGhLuw/z1EmObwmYlrS0BX/iU
NRUvKk6enPD2SwDGc3MEx1wGo6WtIk0g5T5w4K37eGPZfgml0cgmWQfwmDTyWVZe
J+SLwLSsz+Eb3/PAOl91WxZfdntCsvg5I8Fy9y1UveBaYPwyL85pMernox3Lm8mU
PNEM4fbPiEoOhXbKaIufqQCzexXXEaC+an9ReMsSbpSnKJQctfuT6ig2/5w24OoB
MO2dCPnmmuYrDs2Lt/PdaDVgsd5s3fHvyQc03n3OIrUHU8rDMxqW+85o4pdl1aoo
blb7LUMY/69MFfuUbxrKhwQGae3nMv+7RtaR2aL60zw8BL0ytPE1KGe/g68N0KYr
QocNlfiiu5VYl1jROkK+vjIYpd4lM2bE86joY7QKuOqtLwayFvWByArQiB493r6M
hvA7E1dA2AVm3EgrcmByjsTXHMXq56csOyJyWH4EFvCWR42nnzcGbHGvgqffUWqC
CN6qytActL05c1bfsHTb+aXulO8UNOR2pwlBrZrFvMHsZt3iqoUxC9YIr0qGNOV4
dX5iKr9yFfuFSgrQrzpRFXbjM0YBAfxc1xWfCJmFWSMNuBxLugELO0TBfZp8kaOJ
6B2Y+mBm6bwyaRnCjPi+GIeVitllr4j9PHppwHkYhlNa/YQnQ7l0bTHd4CFJUEtM
fKGfBTtZII88DS33ErJmexXKOlszJ6YE00LbYy+JpqwuzD+v6Ul2TfGQ/3mfiQGw
1msW4vJaErrOOEnW5Q01DT5CIWFN3h/1jyKyv6jWCiEpgOYyxGKm/ICuVwKXgnq/
e71rB7h1uM/ZSKmv36hPhO+26iT3J1bVvxqox35F2g2CjYIOgsiuukJ944xtngxa
qQiFDsOs070OUveK2n2AhCEd+LnaE0lrw/LH/fcLwLJCkAgmEDzThT7WBvuG/Gne
kI3ZoaKnawGrSCXVZsxbCjEmegkmkdqiKUGUsVd6rqP8TmmT4hP2DrFkCEr/kzsN
A//a/kWjHsLHrSQYsdonafA1/iwilVnnqx3eOI7DR0g3UTUx8z7wpuF4IPqUiJLJ
6AseMHM2hO1vziCztj8s9jQy6FPyBx06gN4Dc4H3EhCI0rWm5vKF96xBC9R1e4mO
3YZG4leDFeEM8ybt8Mn07V2IKjrQaM/WWYYjjspm8wE9Weq/9t0U7dXy1nrF9/iS
pO1/nwjqM5bdJSUgTuDuh49+oBzdoi1lMQ6FyUTHxkeOke+wsssyt3di77TUvtHi
n3Zc7OuGc0CtVh0lhRKYI6OvaoWPg1fQ3/LsTytIO8eT8zLNcJZf0jlWgB8PKtXi
0Rnnb+p832tiJ1dGe2Yf+jABT29gzIMNEH1a2gK0Xxvlcfe0PjbtHCJhq2lhB2Hl
byuvdlYIlWZvouYrwebG1wC2qtja3YHx3CgpVM1+OyxieuN/gDmLBuVzXf3JgrWM
5Vi2mxnBFPKk5Es/6ApPKLj6iW/BoI8IVJ3mk1z6plwhUf3M3VsGx4sep4oitnkl
iuUfeXbpD58REYoF82/WzZL+u42tvbg/bKVgc8gEk9ploxcskQAQm42333QfQxEc
JDEBGOsfR6Xa1oCjsFSpxhxNj8VARfKL/lahe9YSNATUOV487tP8oMbNATbHoqC5
3C0MSWNf3DhhHGfDkMKGhFaTHBi3j0LYs7J9gF7To+aFYaojyP7Cti4NdrZ5j6HD
mrjUeKaEhEWsUQ0/yM4Wvxgmj2VUWIPd9qCp55pl1Li8EvUbkUI3p9XPCP9lS1Fo
0zAxF7ZKs9ES4ALdWq93W2LpTVjX0Ea5E863xldovPgP4B0fiZ/dbkSL7gb9kPgM
2sDpjz8z4c2yGLoUXvdahqIXSPJh9usJS0yIOdCLQGAKBNy3iFsG4BZMNBPWGH8e
wM8fTXJEXeetMUVJnm8O8a/X5Eak+HKHtcdVWQUPxb3kaLnJZOzQ6UDtcSI9dLSw
T2SlSHBQ9cRjq6EyhSXy6EV72TAnKSDFuT9dI1+w9pgKZFQZa6XpwP0WhQL15ayC
w81Q5gfow0UsfwWvWNvBAUOzj3C79eqlLMt64YomZVOJRLC4wq4yFd0SwZQ62OWi
PVbHtHAFyQJTdhnU2xsFT6o1wdv59BMglIr8eNeeAfzX2aUFQttmXAbE3ukhagAV
NsghqLBMGTk3YL7b3mlHYRnZcl9U3aRjD76P8rs8k/CpHchmebpEwfGrWhYzIAVl
/k6CWIcTB8SHo9ljupM40CjWh02u1kbtYE2puqCPTutUP3Un07Wpx92dONT0OkA5
CqY1fCzo9KZxPWPtbxiHPzcrIQrJ+svtuLjAJkuBGVGw6Q6HdI3xA0iTvqkCIdyt
pxATChQlfLymaUhAe3Doq31QOPTKsqwzxRSTZ/Uf/I4yZVqhU3ywWvyVls3tfdb2
7ELlyWXxRPGtAI3ncA8ZheZTX3ugVOHQn1zGtLGR3deeHhFLDeooucSn61zfWrCR
hCodbrog8gCkD6bJf+bhI2IUiN8agNJ6KD68Hbmfj92oAm10uRjED45ty0UrtM+m
xz3y23A+VyzD7A/67zCP8fftedt6dbk9ExJw+Z4smy2KMQ+4BeW99hkv4wIRcTyr
ZJeDbsscRycid0x5EDZBB45Mw6Gq9n5/7rtGkrCsjSTiJAv/WauXIFsTlpU3uA2X
L/ozx+KoOOm+xVLLk4XIvoaLxfJWWmaW8fTB7IR4il+nxxpGB81zbjx+7PLsH4pb
SPLD9vvzIyFfBj7YJIsAklw/8VVoLj4HsFcvV3EiMJnz/A5RmRPSM2QZy1dAsbem
euK1C/sTmEVj/oFUhBxZg8c1fH7REVvuWDQySLprQfFVtU/YSxOJR7bjOCVVdwXJ
XsqAVWVoVCH/VsgGSg0UXuJJ0u0C0xm7+znkBYfyhntQZa8+yWgDpMzgCE+wyY0o
+BCpYJ01on9pmBf7rOrnZqohHMKi9MWnuQwBRbfnd/fTX+dIIwtmFod1sWrZoku/
XVz/+JyDcI0GslgWJYmWU+bor4VrIcWtJ3sZAyAkj3k+UPSyP0TWjkDsl6Q6SG/O
AL1OOQiJOWO9cxVsMEoh9NlJdrFmZv3wVkwD1FJqI1Bb6ZYEVb2H7KyZWZAVN7vf
NQV+5Jd3IqS8DSFKDr7b0Q+D4wE9aZtJ6kuqRAtKsOQWtWdt2A1lehr6Xkc9vqGW
azp5fDVe1bOV/xeq7zr5vAlntTo821ZYLh1Yurcj5NxOfa03GDNWRa88i8KL9vuV
PNEzOemAklRKD66GMN+/njSOxJFTHlWheltkxkgidpE7fPOxHvPRKph/KkyE7p+5
dV4bexQmbWq9D2xU9BNA2JGiT4bhqMwg+eBndvnR07WkSJ3QF/n9JTnwXsrz12hV
cmB1ksDj9GfCRNL4FoJfBicVw8ktC1lR+2vP9hwOohXHJqKZuazX0we1tCXZHGsv
S0H0hE7l2R4yvxdxn1sWXITDP9JoBh/nvRtL6HISILSZk9mi3zeE3Tz3rX1RAFdD
9Xog12ca+ZVNRi35FondxoQfpnAI2CO9Ti/H06ikbI/rMXyvHDRhRFlr2RVjO5Vm
VbUKKAlzMGXnyURWiXIhD8FTMuKO/7JqSNyr7cxBaKaOZtrSsE8/sMo0yDNsLJPt
mbyGBaJcQaKStCqHRoSlk+a6mSgnm7PSN+s0vErx3xyAYo3RACB6CCpjfrtNQmZm
srM+25N/yTLDJjYKSJPV6r5bMp3x/NiwJ1kQKIavv54XOJLedFZwG+CDj8dtllmY
/oYd3sH9if5hYpTDE00B7/hi37q39dvDUjH615QmPGf2gXdc+q+7jl7SilY/Ecbp
YDcT/ux2ndxB0CMEzPHh3Fb/I05EZ4JvdwT6rFFzxA61jj/qUr5WPQ6NxnT968gI
1v1oM/7LDuwbQdNTs7XDXdoh8WrMTg+uy0NjxcCWbbq5V1437O6qCCOxHBgD31D+
EIHZ9mbM2g+SCg8ibAZnRk1VClDS7udmUJnytcnJ7sEcB5+gfrfpz+mUDLftAlkn
6dbA7+8iU5V9LO0Q+fZxMXBuXCSb+fOwmiY6nb/bLryJwoeKya9iDC1D3AYgNxKA
vU2aCROf+us+zspl7vRhTSJSBxavaQNznJk0CY0A4oDEkj4kbS2Re7ICFQYmh/5c
qd1Ioe3SxKZWf97Cc0PGdYEMdRAjo+SBN59CQA6lOrVBkiJokUqkOSJ+asN6IbiB
JGNcmYKaGsMNM9VrHZgd3+77LgTKxvMzjauDgKdOF7Sh9Mmplr3/XsPOe3UHm7yl
XD0whaaLRxb1KI89CU5l4JLX+yqj64dgktcqg2i05lwcojpuzG/VUsradKqFAHH4
3ORSORPHW1GEj1ndXfUhVdB4H+PfG2ETMBG6Njs+65VnvDoGfxcFVoHNBKrfOKvM
aOmJmL0Wa1c4bq1/REbJ876PcmE1t2NgrcoIZ3NXENHm07Gl9uZwy5CBZYFb/+2j
QxKg6cyKX8j4kbXjQM5UU2bMk0M8l3c+tdfKlcs8FUQRgkYpNvM0nSRYfVuHwl1j
w0wWt3y9KDlkzoeaylIkTbKhYGzpFtRC/6waWkSjN7zCUn7XKTmgr79Nn5LZMtch
HgsKX2eTaGjPhw+7SoHWmWClPA/QAdHq2X/apGvnzTw907FSQ0oF9YZhJ3Zs/Zvx
FxBfk206flh2uxM0uY86O/HdKyK/UzAG7s7L4WOlVy6Q5oAO0q0GFNHRz3qQo28A
Cc1OBYt25+IXT+OQ+NjawYspZoc0KCtt/DS7kDTZqha1Y06LMmaXvQBkg34/2msL
P6H4dnJJopQoul19zlBGut52S25QTtJDCgFVz7dgk3IKTLnfPwboQSvD+GSXfT7T
YA5w5O5WMI8snxdaoZ3l7gJROrji93uYFHHiaL7TCqykzG0LpuE/Ss9rV8WlljGK
QgxfcoyAX3fVk30ooJp6pxVRzgLGaH7V0dUnhTGyCFfje6oDENL4hmZLY1/wTCtl
d/Q7VoSL3okuuDkbgSKahqpPczcHxCd0Tf4ldqr1FYfRtCPAHW+JBzodYHJFtTLX
9ZIy6A0SvPuZn/hTr5vSXLbozyF4UQ0mPRnFUb/Hlswc1BVO80S9kuMn1EuCQAMB
zignZ0ToV8/2mlSO7Ho4O11r0CAaz5dkW9oAanb550tWtus9kU3J5thcEYDeKcmc
NqzwThEc3Jtoj4hYScc+otUpA547MeVn46K8mgjx5q/fNZpjVZR9augiaG8RjoO+
07rs5rDCzPpRnbrAdL1lobQC4Fu4OZj1L3BY72gOQOkGyOlMWFMRlFZLa9VSDa3Y
C0Sft8W7ZhdurhJpalf/knMIRNSc5gUVOuu9xitQsUElwYQdoQupaLih7kTdoCDZ
o4u29MwI7V2Z2yf/KR6bV/OaxWZzUiIAzb0/NwWN5xA7dzTLh2eYFSLvPSumJHaV
GSTVGAaGuYkZVQ7QVZcdBYiB3H3Q8ZkHAL+Nd/v16SebI+aevaDnSOeL9yyoSxDy
k+Jaq/j+J2e/Ychr4klbpjCrVj4ToVDs/KdIVtcDoQiHYkw8DzoXIOZvqimz+GUN
JbJZvUl1JH640IgXfyi31cc/wBBqt4n2AiLrduqogCK+Te8sbInJ2zIpHd9I5KN9
mh5Jo84CT3kdfukBZ8Y1sByi9D95HssCOUcBItEV2d7zfgSvQ/3h2X4yt+QJyv0X
vNXqEVFhDaBD6cxuMGk3W54danKPQNcoCmJVg+8rNwqKPc+A9XO0fTNvCNRNkdpH
goa+B9wd719BO9mZwGkohPkkvNI6oDcc9oOwefOP90e063h185a43ztbqka1Q6Kf
uNHnb86s6Qpx5nUwLX150EgHkl3IgBr/veH4JYViycA9HUYVd++6y8CHTKO4ayD3
G0+kNUahEo7h9Q6pcwK0fzTnUvO+KUKWPqxrst1nIBZ1AcWtit5m7dx7yG7dyZ4n
2IrRTYQIDOqRGfRG0pVlA0f6fASJ6FT+qFdCV59WCzxH4dr8O83FJgt0YeVfmhWR
K/JLUI7NbxUHbPu6Ba1mFwE+rBExmbY0ZgjRB0Sych40hzrGLFkLjyIPOihyw+8p
kaDXB6BjARIPqbd7lhZobJFZps1j3kffLar/Ow1lDpne5orJE9YImPbx8Qvl8leC
KEU/gKw9DisS1eLVVa50WH0oVyBZh9PJMraTY2c25ApIeAIR1rm/ozVkAtcVEuRU
i1UCd9puZPKCIJ6aacFnkClj58V1YrIbQfaa2I2Pt67/Z/Lyl001b5UlE/z2FLMY
v1w42eo/qrAwmvrmUwjg5XHVMLsrUegEagig7ytS1icCU5KEgl145fQUGknH7n8u
Ttb6HBxUhINQ/xjBvReExpzYaz7P17BWcoYTykdW4NrKFrXEmyXf2vfqNcoV0vi8
aQCFSea6WA03+tJHW43DE0C17MTkl9V3LhmM7HBD3tl9BHeYwRc9tlkz9DYUogZZ
Vb9PDcloeuk0Yif4zPxf8NY53xIjke0jxr6VWUXte0P+/zBJt5Nhir9foqBtNwS3
oNc9KSEFlDyUc5Dv8Y04isZzttL+BmUnc5umQsJr7mIZ0wm3CCeYOG5u6H6+B5jP
dS3ePKAYa4pWxoBqmxoLENmAGUkUuAHYCC6qtNsKN8HsJ371efvLQ8+PBk+4CYmo
YX5BzNrNfKxeoqo56SV+VLgc2S2TuLZDV1ADjaZ4wL1NC6XhBvn6ZGyVqoM3S/Lr
YjPi30O8d04KgPIihmIBlIQdMUHO0g8EMcLpvQ5dZ2J4BQ28uYUfuXVW58CFY81G
FXmitlfPHcVFYNYheYXxPGVLq7bZWrMAEbXJoNYqiqWuG9FWqDrND+KJL5qff/yx
gctHoUm11GH3JVsWy+j9X0WFyNFGGaCUPuQXA+t4Z37ZY5vRJ/VnrAoI9whnPlfq
RNr1YYUmzpyUwCQHireZWzN182wjDgG1n0+Ysc37y5sKgAcFo5luzz+GYh6x4xq6
NJUP8O9rNMzfZXaLSXTeOe5s5BgvacrthHwca1Goh3qWbL0kFQFttz+FNHsNihKY
2W/rGW3QdDzaKl1WZwWPVrF3klQPhYh6Dv6k22nTKAS/FA8PUZAADZvUNANN8G23
FWwjTI0+svWLppaX7YoCewvbOek7krWQtcRcZKS8h0YERZS+menOTO2EQclG7nrJ
yJD9HsExGesH+oCw3mrwLD6FUfLsCldRwrK4TE3J+ZLDBaXYNo6GpLj47+OwSBla
9JSXf71gqtsGo28mF3h2Ao5V8CR0WxgaqzcoLBeQuN7e22nAXFBic2arEEFgYVVO
sYJZz5PIcvAwTAeSdSXVyMgqljE6CEn/ve1nnSqVoSp+ox8/t6plqa1C71RmxNcn
rBJMEGGboCAFxtoc7ccXUy0/1sEz1/eEuzNrRFxA4muU5RpbX8JOWvSVqMcqxV/h
khB43q4FifWr6wCD1cPBVwfSNw+lURBgqe/c2Zj+qAqUsijoIuo4BbNQxNj8py2+
881EoZ/A/mMcbFRZT+3oEOhsEIoSPVSGL4MrxkQMmpPKX3Xxk32i0hi2EtW7fdeS
/Oz3DRXdMIW34zp9tjc83kjus6TGyvFRefIbJ4ZqDiE/gCOOn4lyV0cI5vfZUV/2
akg6gUbrsuwA4clgvGpGzojNfj/0gg0ZGzX7mAS6Al3bGtgglj7H7GY9jwDQc7A6
5Xl8lR/P5ncbWaVU1/d8v6fChRYR3Nkzj9PZ5sTUbDM7tO+a3axUPwg+vxy4oqCf
Uf5j6lcgFDg91NL00HoPI+hka1vbSiMr9bigiV57Xm+fWa9VeIAWAVpolEWieAY8
Skm0/rwZk8DT+G5FUbctIJ4TGAovsmHQcQH3q2KaZLhuLfjZGyEi9+IrHaR8kQHW
bv98L5TAm00YZg03TA1wLkD6VuCPe8u7qHn5In35AxAU+QVVrv2w9QTCOpWZ+htc
2w1jmd3V6Yyh/oS+XuW9T1hxQgunPIhvoKvNJpzVA4hi62zUa6LGelsAkF9KbAsv
lJouRX/FxqiXFVTZKIig9vCfcFGV3HAPEmLoL+vFRWkdB4uGw8buBk/PeAt50MWT
8WpMW22scPWvDJNZ0XlYgRu73M8azHvC3rJQiY5inK+9+rm39VUzpjfbXa6G98mZ
tRzzHzWYgTcWo/bA8lQhxjk4nvO37U+KP9WKqce3xhsJWnoxcKZSIkEEaAK9HTu6
/yHdRe+LqhdipDFjjPxtiTbnliXWAuBn0f0yqorly06VlZduLKtqcaIFoefXXNGv
3DlhZ/LYuNGCgbXKav0rgIC6HeLUM4fw+ww388feVrcK/pgRN2Q2sqpV8nL+MVU3
NzdV5/4y6GyNuLn64XJCmFnNFh199I5HYOBJBppVa53DIO8D1p9b+HW2UjHtSM1I
u6ggG5R6tQxNm9FP+tDY6kGW79QvsSDzo3STzzOfH6THowWCpL3DVVvVwZr7Ob0q
bBR9ETmjNezxeWjjzuIv7m9fhjKXw9gypxDA2pWs3wWlAkkzBGwzMflJDmDK4fMx
+CNUx7QfRWj7jTz/2L/wVA1gytK5Sz05C3u0j/TA9wq5+hFhSqvGA4NI75WeIKNY
ZkYDTPL5/VvKRlorrlQcLX+ODmm3BgFSg5QKga3N35vY7WuJpgO9MAtEH8gaDrf1
poHN/za/JLwjDwMZ+h4v07duujkcJVXFesKo66DvRnTN2JNq6Clkr2DXjjkWlKZx
UVMtNwQ41V5y4xhHrOhKDspM17D0Kk8HUTkXHGoA7HFO359BqYYBuo1MtZrJ6zD4
Ks+w9028UU5ZqSQYuMGNUROG3UNbAezU+4CbCXg3z8RbTZItkqlhDDULjCgqCE+O
W9ggXbDShRfdbqlEShJ4NDt3stu43bVgOR4E2If2hfq2mPW1oONe4+sfE6MFbn5n
ZG/Qd9vn3MAhw6yBPbk05GtV1lFGaE9eItm0mtxk/OkWHczhKI8XhmyOSXUbpQXe
DwZsxtVxenJAPoQk/WcH/n2ceugY7FEea6aYRRHb7/5nY/JVnALj7p0a3z4YQXE5
XkuxG92eYWyARsUKh6ormAfut0Lc0X5c1vevr1O0yj7eGrdNfbX07l1EcCnDNW8i
Wwqwt8kHd7U4VKyFz4S/Dzxw9IF9A1BfhUggCo5L/bQxmZ6dfoYGGA0YBKAcZAN9
4ioTvcWFTaHbTFogVw/dVRx0SfrMXlDwCdsoHxX8iowxNhvL7meMl8ZqvHHJcZYA
EgHiVA8p8cVligWjgshTK8EO7OBgif+iY303IrKwMyUb0xUfJlLOgJSlrObToIOH
x9YdNWf6CD78WQCBDYRqMNZWaB/NLknGcDk3iWHsnCMaPmYJgEoWqu1esEMXg39n
0fZNdK1tS1p+fO0RcG0i02HmnPxI+DMFcyRbbGA3Vnn1AcAS2ARMOcxzHod4SzSZ
RGVq0uTge+o1PBC33hWS9Hmy0JpYU8+k5iojNnr6qAifyqAH6jz+SUPgqE159sCU
36vUWGiwtT6s7AQ12zPvoV5xzLCgoqbZpfuFGou3jr2ixoKmNgfDP7HkRsfCgggm
31+gB/q6PKbw6bemwM32DRPFP2cQOGkOJszlcUbsfkl+MMjKnPrRM3KNy97M011t
hz/N8PZhIOlAHv5CiZmZmC6+wulGNC7mDYR3pnIMRdd8k18Cj5ayU8Pa+oTQhkLi
yQsHkbqQPB1s8bjTRYBO4BajgDeEY7QGtYPitc8Axg9UcFWSewLCu/frbcXozmpD
884AB3YXMtuH91Kp8PgzmhtlkAEVpGKnYCggFR/71iPj8pziHwob8YJ8kXKLfgvu
oCFppLHlJ0ioUt+Ct9jmU+YkY7DjcQsob6h+bux7/ZqsVMXP8G39Vjl3HLFxJKgW
m0bfoUFI5EH0+KNya3YLzOl1PcspxE/RExnnIShOSjb1cD0gFRliRtCUQ84B4u+w
FisZma2cm30RQkcIv1Xh/Q3A3uoEF6ivo2u9WbI/zt0lKaJWubmiU9mw3aO0EhmH
IQILSZz5XjCQ7UgkeLGgi3/Yq4G52J5NpFF6xEFgLe4zPlICTD4V0xIY0U0Zw6dv
KYM7SuPJLFE7fNEhkeWh8pcwc0kLS0ProXQMlWR6PTnkEabIVaI2ileMUgjOFYR9
U7sSVDElJuZ8p+6Pzf3Y8jJRrzaNhK2IAKMn8cF1/WVjN/FIkd1VR42irpV/J4uQ
riabnmFQnrgNXmH/muqHvoTtT0xqdyxNNdAS3S2JTW2DtuO5htaPdNr+2SiOOxSR
tOb2y0wZNW+WRpxG3+fTf85ZE3XOdGW7GBlaTcmDfyv4gDM6hswkRC3odvnKHj0E
EtGhcVLhz6/Q3ApiT1NEf1/feMi7ayK0HK0wy6j44wilwPUT3wlSFYoBJNQDe5wM
By2f9V4yXXwHhDiw1nmzwUs8SBOyQ1xuaOBOSBYgBVBemVcnbOBuzeLuOFm0PJvc
OfKtOzvKblOF9aYBNVKDZYfHjxdPWz/NusdQTMKExJxQKl4SL7EH1pEwcJ/VWKJK
mZtpRmPHpCNXr9oYa/JAQe1j+m4w+bnOoGhrE0VXtpkfRT6T9lW0rlUVuzYE9m39
fwuQmkCsdO/xDi3WwK2bEiJBCabHxLrEv92pf4TOy5aJ9u/CqxPmxu48kEwEBdq4
whhC1Ud4EEVbC99CZX4vrOq0Y5dp0cDJYxBVUFeWobf1uiMSi2DVg/1m9fuEkH66
i2I5BjHa1HTA2Nt3s6uVQNl8cRByWsVxIbK911xDVBPZr34slk8tX2dHiSwg605E
NR3KlLGrvJe3KWOgKntQPvAf1671vsh/YdNzeSQh2ieoO6JhYmChXl0vD7EidogS
ecdiV67KpfSiIwv8SSU3gI3u6r7SyP9M/cdC1lJeYcvC0HLG+3xSJhZTBi0VRI4Y
yN+KEaLHysA5SjZUjGDmzs91IbE51+bhXYzkIjJGFQIewiUhsPvdSoBSBRl0MtVc
j/cxuJf+SYbNdWo4hQf4j0ChayOvFQ8k+nec69l8dhpZDt517zD3lLwJ4MUBjMj2
oxnnFgIhg+tZQSMhy2VJbGiN88DJUKewbXB9sANplDshyRPT+dY5bh8lO1YUwiQ+
iH5/sZprkEWtqTxg9rsItV0yygJnkYBlvhG4mGoAn+jQCmHQ8Pz4xI93R18/f0Lb
CGPtA/wgFcJXM5M9PjYzaVBv6P3D6YoKvqYnQw+JhH6PmxWgROogdcPetxSa2jN4
2+H7yEmreZ5VTChVR9PA8k+xQ67i5UoCyIcx5XHPaK6MRFjOLLHLYQDKqhwEpJbv
5N/sxUljEIIsEQKoYxRK2u2e3T6l0LwBkOejdreKVjN4CxO0WefNfIjY6AuHD+Ed
jBlp9DZZkZF+CsgTqnVIlldIFvTCol9m5fYlV+DMa6oBkCvMRSKKXHS/t84wZNoR
bK+2kUdApfWwm4tUCL7FQFarDWxtC71hjMmtb/kKlvOCUfJ/9tIF8xGgT+eT0Rog
LG9CN1/JyuKoyeKc+QTGDE7Pm6kp0kkN2Iq+RjuEhWjnM6fedNuRq68ce2SUwpta
LT/95bog5BjgiFOaOD3isxA1uIkOkbmaNJBZrK8eTSI8dk7URScrXRJEiIEK9rLG
jx5UdBKKkXjHKYDvQ0rv2mQ085ocFe3YeuRKCE+kk2xNYP4j2dWJ8C878vOTI7xW
B+nhsNaLgTL7vKCIyd87n4P0fl1KqTFBnudY89Ss0bnydDopFeVYpfLPxqVqTxE7
xRKI8W3HHHttAvdtJeJs46Jb2BXwPuEoMCptsTCH5/bM7fME85qonVh/pcvWUNyq
FsA8kzK9LzhgsIK+LS6Yf57wWJDdpiSTNW2CWPZ2UvO7/wldNqdBZ1qbYsG6DKCz
8m/hVg/79xf2RQ9/UYbzFyHyc5VMkpRQQqeg4n75LzFxmp9TDJ/C+AWYV5LUGFei
JS+TAbCaio3aUgHt3q9TDo1ACIET2lkGOXTdlsFXvaFzV1dfuIqjY82YrgGwKbho
OT3y18znrE+o0plqeNEw7AXhAK0YEtg+7flufeg2QnvCeLsjmLQYcJSOE20CYxnJ
AuCYNKNye/6/xOb3mz331wCmHXrK4QrCcDL/L8mlDeS9lZqUMxNYxFeNBBkVfs/E
/D2TRulwaz8r4OeTtUfxgiIDIkdOLTn4M98Pfah+hr92pyy/uNbcSKH79CeVySRx
Py4y8XtzJFA2eLEBYstC2RYXQNT2ax9EqLAHcSDEFjYERFZlO+D6K5mH3Air7aWw
a+jwYc3CCI5Knp3t5nlKHCgbIJ6zbM4EcBFgJv75Tf3JoKxEn3KA5Apd+m8Nub8t
vwLv2CVfkCJBqPwrem+YslBDRQYgnjAo75URk1MfglcHWMGWkNJxWPdpW6wjf31D
fTyAHKngyfx19zRppTwmTSjhJkxktSM/s6281FIANYTmg2MlgU4WUHG+IEwm07Am
K5hinuWG6724e1SKMkDBJSTvEZ8sRh6YYxI7hHAqnL7N48K75ve+BRDGzOiWB9y3
R0E3qwDMOcsFDi4JQg+ZUVYHJVzoCUsLjfimWV7k9cO7uIc8PJkm/Piz7LcFhIg3
UaaY25hTAp7/FJHJRoYpC3S52Vm40+hV72d/u8JYmvEAlD334H0MgTXHYODfTLzI
3NHS67kQTscFMVi1uSNli6q5VAAj41QtJd9tN3aEOXLfyyCkyUTbLRCp4u7OXpnX
1Y1WARj7pmLYfTq3kc/jT1hYfo9rLTpKUfU9lW7NvvP0nYBKMX6H+xz6H3JF8U+/
39VAhgikzcYEoDf7UzCHXiL6yaN5VdRMFaw/Wt1wlpw/UmGkJ3vmzAff/iw0+Qfj
Ws9cg4ayzPt6aMk3UB2A3+9PTdcvDDHw7z6K4xrmSJ0F9M3ekAfJWCaudSfXInBg
BgO5mZSNUiDc9T6xGT4GiaVfcqG+uN3JsLz9Nt/6q5qmrHJG/VkMrcn/gfkErIN7
25IMV6oSB0twBILTKuIVyYtxdjK69I30ot3fQxdub9sOJ5mTcdOCnZYdvRy8XN65
6lkV8kglTxd/wpYN1H/08a8xIMN8o0YN6xX8CZ+cHprUumhWEcv+LRrvGvTTmRIo
Rk5NWWqiUIUhHUphVW6ORkJts/vCQtS2eKeZ7ychtqS9CZyu1X5RGDZwF8uVCfpb
smPV6u2/cMyVb1Ad5blgtg2sGJuqBdSe2HAl/ajyQpX0+0GyC/kE74k16rJpG08V
byYq66SaPSy6d31PdqgoyXfwH79CPu0NDF+B6PieAajr9HJs+ATGFfX6ULlGm0Q3
anCwGP7OROnRUwvnfR0j5npoSyX3wy38DdR32GNnqhQexsvOWJ0HCY/GzqyK/QIt
6g7Y50ssHGufomtrvYtDnck3LWXSHlH5STADbm1lxmbeujv4gUzeVkYjzb9vxyuY
6/UowG2gEYdgF0yY58taLkPuOOr/ODWcAvPT68t0T/cNA+YdVp9k5nRK9+0hZuhO
7F4+NjExtMPhW3U8V6+w/ecSYYkTkADEfzdy1rHNz+TmgT6FmkNzaiEfCok21C8a
oFUdwDcJcElIlWc1feOXDlIvioCU+QR1xP9F1JnrUaiQ/GS6jBPuaERCJnqjKKYJ
sGdnnNKLuLgIfpelw9jmteKWYFO5kqZeG4scprBua/eIHuZcNqIom4yeE2i7OjO4
pcZeTTtib8ALKtQV/ldaTuuAhA/DVpO00JnG876Dck9SXeySYYKw9+JWNxAebV3J
UHWvtBraZivVQQrbVu0sYtiGuRsoEcXOcjk8Ie4Gv1idOhwp06YOF8awOhQPspyp
c9rHBCgOfq+7OlhMRmYYv8NmKsqCxK3OakGbPNMh9nZDczOv6Qp4ygDV+f7cnvu8
2Cu0XmpQ3gWvJ9YO09T1ABNwr7yMhc8H1aPY7iCqfa9ccwadDbQJFJolkcdmutlY
gxCxAEpn85STN2QChszCk7hAH662jUvWZ4tXpQstZjA1OrojNEzS7GHUX6Yp7dSi
GnUZF5VW5tXzeNVJDZ4fWZWkC2dBbZnrcx9BRpUgL+zgwAhXyYzBRSz+t+GXxfhk
VYpmG+ya1kls1Vc7EK9xjzDKYlluEPMvaloWi/i+QjLtubckC6iRL1knZB35ppKV
/QohZCr/VVdcJYsWaBiFiYOLNYuIhh4VZ51ZnV9gq3G+cEz0dJLw+6M7u4FMhSZC
U0AO3f8V0VwXaiI/OcnVA0GcqqNn2D6P5EIGCZhUNSGa1XqE/gbOyqqjrj2mH+fr
rUUry9SB92iZ8if4lodr0h6/7nTKSTOQQsSN/PEjdTH5PNzdXmU6aSkfjwmILBTv
3/2DBzmVKi8IKZnkm63D2gx7lr5EdrsZoiOaJRCqFx68pu/eTfa0gg4X1bJnsdAk
ty/x7nSmOTCc6oIMO9WMDY1cC3PkOSqjJ06C2CsqTAGRewvKsCzKW6CAiqxXlmxt
09h4Nr/dqEpugCarpXbCI/SMtt6AqKjeLoIX+QalX+b7nh5uVs4ohMLRwehRid1u
1gqBZ6Q4MivDmLd4ruRYSLoyP3/JCdz0lkI0Q6ghxYwn9xNWxVu8iLI8XnNF2Apc
9kFEqUbPHESCI6T15OhzpnRfrdX+c90hZbIBVc5zEU/vybfBk/Nhxoc0xglEjztu
4VTBWm62wIo1eEcHF+Qkjodw/bjqlzaRmsHd+jdeLfGlNw4t1ArwnTGZLswEi8zN
FLKW9Dj/f5Gv1v0SI7wjFeahDLxnQXAPxMMnNklVrXR2DIemeTFAvBDanUmWGLHv
uN9osMqVBvtGUSNrmKl2QVz3MIQ/g2T7vErTOvGX14mN+RdHTiaw6bsmZOBcfqTA
sM+BtKwVlC00/T+viiy0NOD6E5iOchMrkNoQEjaNrE5JGeAcsX0Xm7n18J7qDluO
2IrU5EncSbX+3KjRIPZ1kq/eU0XsodwLGH7nV5yS+5rm0CwNAoS/JTfR5n0Mm7P3
EojSLSrBOGqjB7gX//3JN3wgxoKYeAUdyHUFAjaSzY7UPGzXwR8QWmpivWiYzpGy
YqomwLe46zs/hwOIBs2zYp1+22m4+By+koy6V7pACCfGyF00MfZGmkG+n1Pz6r6n
JcTqxeFafsMLGO/1VI/Ss2zknI6nJ5FZotjzwY45QWXFrZ+ItPZcQYfhTRsc1uPy
MiFYGSjcZTuRV3mnCUNNZE3rcE5nb+ChO4v49ygQ51HhXgkTsP09kXiCuum+L1fJ
W2lZIVSXdbaKuG+Kt8HrKisFQagSN5bosBxvEpeubmr+10u7sQbn4ZzU6QUurZtQ
XPYrxvxoSigVvS/RbIBRLTE3WCSR85bSu+LMRTkr09bMY93v74tLSF+XpNvRc0j3
FSR7lY2+udiZ+RHaLM3QeLlSbHYCKlDs0aa1rCmFJPrdRgQw/A71eBAwUC++I//P
as1IvngFsJ4fSK/g3+Hv50H2/I4BQ4LjrUXs+TeWWWudLEPNRt8mnk09dXS5mkPT
AOonVUfqOSQxNtf+WnCYNH9xT0VEQQV7TphUB2LyVa+11C6a+5IhLUIa12IyD694
LhkDHTXAVuX5HFlYN2d5zb9jFmmtfC9KqbcBl+C41PT2T7Gt6F4BuKpsq6Lfqmo+
eQopZioC4k7D7iRAGJcGWtYIiAe2pdAIqvy3XMFxcc1Y0/TO7YaoMbHOu70A1zdR
HjbU4Ucdy/M3Lbr7x0EczM5Gsr6QPB6bdp7SG40nEN8o8pS0eHaEPqapkannvXzK
wvmGbxxZvErInMVRSo5wX/mtVs7JfcJ6PPN2j7TQFQmjioZuK8LzOxPQAWwRjXKi
QbdWb5DI6vQk2h70RWmeo8P8ZHTuvPZW7UmkP7RQXr5jBFwFRE4FAfVP03IoYMT6
J/ilgZK3I0cPIjqBsBYbAmIgIvEAl/FlLNHJbA9n+76fA/GrXedptBUsEFq4BMRV
zLWsJ/9sVL16pNT+zio00md4VCGR9C6ScEzacxNpGCg+IEIsApyuGmewc2woJLgm
H4Ucq5amyO9hLZq1MJ1wHkwM9T02KkeUkj/JxANvn5gIajyqswCnKAy9OFhIAwQn
6uq5SGFH1KghGkfk2X9b2U70/Vax5/S7qkGgwoESPVc5r5QyadV+lJledu7cAoAi
ibPpqt/3YCuTvIZNZHT8O3lE53XJtDynOl6bd4SS6GMa85pasqUFX4BRPJZclP3Y
kZXdf6G8q9KMwGIBKP5NYZY0cAqNjAcwO/qMAo5Zd9GUGyAPhMitMKsm6qD9ajZp
4jSRTzR8MaVZpZo6I5ljKS4oSfa4EqVJ6Jq6MeViG/FLMRvM4knKpiClwDeJMhVy
VuLRtKXbNLT/fV2IN9nUlNMtZ96f85bl6zUi2LidkOjENBQacSllLL3UJzRN8WP/
SJjmt3pZyNWDPEQv4p6CpW4QIQis7YFdeJLjE+YWqOrcx3vgDPS0reWFdRDpwvvd
3VyBooPL+ipmb2OBgmj2L+piAsXSHgpg1jaK5IyPxSa7PRXJu02L/WwuXV0TTdIw
4lf4s4p24eqwdyYgnYnGmhZh6TUqgqtyvSSZgeeo0bYso1Rk4VswyCwJ/nkyEmAF
BaD/xtCvfHjVyHwvjyveWDWN5ecwtjdJY0mEEZiVfh24K21+BavVt4+DDBRJNwLa
FaEGw5e8lJNEeCqLd05S5aKhe2gXqkB2RRJtLTUmxaxD4foVNfvqelTCnGiY5hht
AZYBvUaEuYxgUvWOCaGzAwPa/cmirX38Z794MRXlhoQfeqoNnHjWNkCUiJpnLaqZ
wLZBmjiw27CbLO+Vue/XH/Q9JL6G4ThfE6EvTz9lSMYO9Pth0bfUIWXXA8VylB0Y
j68dricW9sWUcXBAW9pH8vTMHWlTyinGpolUoIzhZvdqAKsp93HOoF2EyGrFiv1C
KJc0GhhxJeGP8/9fhebx0MsDekfoglBU5f/0Z232LRKs+j3PtWsqFJgFfuKJvTvi
OBYzByC42mkmEGpQMlGocN9m3erqLMFSjZqec+JZUFDzgWxUdN7Nsli1FvciqsAB
qUkpyNyNM9yt2+pavNItl+1ySUkJmV2MhKWUrrWSjKttbZgB5dsWDMgY+laMCBzU
csBRMSz9ai1a1NJWjqzJ711jf+FuKqS9cTCwAv8Cq0LBupxPjwAVYmGrupBCMj7H
d5dZsZfv+9k3ev6Vwxap7aR8+OOC8+6JOqnoAzWE1BOV8Pm1wPNVefvkEmNbLHGf
BDqMbkIVSgZCJvbq/RVrcMnDO/AT9yqFIG5VfGhmBBDovSfMJ2qMvBQ9k+GgynH1
Zj8FBBD+3Rkgku1hLU3f5jqXJSi/t0LP4zBsEugpSJ9kl7em5yOlAqNVrawpRmo9
aULvOQVqOr/YNKDkuYpGmp9hiEEBSHQuaiXfGNHtYpcL89oFEXzeFGxw91Vth5CK
gomh/uUCACpTNgFhWdgk6PWI2iLTTY0ODiWRur229eyBIRFF+XPnens+brMLY2tt
ySR0SUWN8NVCXJiKHhsZ0diMi4pGMu/soOczhW6ArylR/OFXSO9ExWddaUz6LGDB
z18/Ob6/ak8tTmRpJZU3FmuDDGm3sOtWA1RTSRz2fc93zOLf5/yjt8fNDcV2/qju
encjnIhMsDCmatTIOGvOaVprNNz0dCu3s7cPnTarC8EOiTrMOPQpEEeAC+4sZKjU
mbcES3U2dapPMGdNwhW586ewrU5FvucYl80B4hvlBI1ROiu8YvMqyJGEYlrR5qqW
TjyhfSqAXfip4WdSsu+LMQyQIMoaHWdgxIvAD3NA8Jk=
//pragma protect end_data_block
//pragma protect digest_block
utCbZHrDpRZyZZSMPBK9wUEW+jM=
//pragma protect end_digest_block
//pragma protect end_protected
