//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5W/jOetEGSXJiBpm0lBTygdvwIuyspbQ7kBCmpo5RUMnhsHPuTJzdZTUmkhDTbhu
1DFygolaPkH4krkYEiMd6MRkroRdczVPRR7sRBHDCIJeBNcLyLBpCk9SOAJQoH58
fn/bDMu8FYsGQS8hucGQuWragEc5Xa+aWor+3UdkUnRqez2N75oB9g==
//pragma protect end_key_block
//pragma protect digest_block
C5cT4Nw/AQlCSOdS4XeDMUBkbXo=
//pragma protect end_digest_block
//pragma protect data_block
TZbdSq3HG8quLLcSwWppOazAOe9uxG5FyV0EbtVlENkZoP46WQwdiLVV1xuhQ5H4
yZwkWa+f50FcprLwwxgGVJrYX3WRL6Pjxe4lL7hUGyxVvZYMt5WprbY8MBP1/QgT
ctHlFfSPQB2dQFTy7cepSLAxCWgPXm0xMdmQ+XgoyDmtv+7D7U0rWJNO/y8fYwgz
BhsJ01Cvvqnz+zaMqG+T3YX+RdCk+Fz4nx+oBj6wGKaDXiKByrHa/9JoMWT5pOQZ
em2rnnq4dUn63Ba4I0SqUR4vcmlgmvlG/4i2cq4bpYoskQgW6hkzhxhsJ3vz72aq
OVNyOADvrfiF47JlNvPOvg==
//pragma protect end_data_block
//pragma protect digest_block
YvGdZYK/ujD3GGiFgk3hDrPoZuM=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7g9W+tBDp0AstURKJtE6bFY+KU9SGswmR80ZRfI8SLQBar3Lp7gA2L077Rbe9hZv
XUee1kGzYOmZqUH+672dknTL4D4m03V49+9bi5QdiEBdrr0c9orqlR2VBpPB1lgt
IRZgrkJxNst0yJ3PMdCP/tOZhfhoLKTo9DEOhmVZEV1yPjRy9wOzag==
//pragma protect end_key_block
//pragma protect digest_block
qyQpgdW1nz5PJxdzCdF3nEUcB04=
//pragma protect end_digest_block
//pragma protect data_block
iFEriLSWqP+pL+Sqx1B7AWptpripzwIC9SE4dKKACGT29xs++rJ48g6Wnc7sf7V6
LBOaK3B6dyOp9li0UJ95g+MOa7x2A4lGzMX5FrriXX3B0K45q32t33B3NV9UhmG+
JqdOEJioeEHmukT5ACq7b+Y0y5p5oXWdp62BUiopxb1PyYK9JdQAnqtjZfrXFC//
TqFhgRy5+t4xfDzpzTBqRNGJIQ5G/VPU3ZQagDPjRz/SpZ9MydyZLIKufmmUCkNR
FB5zI7HZ0XCaSGjvee4zV++9c+0UszzGxVMhWdlQ3d8glG1Bfxv4CCox8vCJZLr/
xv3s8vFGQfpSbKqfdeZ57g==
//pragma protect end_data_block
//pragma protect digest_block
HxRXC+yijjwyIUnCqT/5b0jfX6s=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
4w/vISvz53FsBycuaH24Ubg+cBSjlX3qk9NCCOk2tJc4fRMYsOAu7otbStSDp6AZ
u8/wd/5i1kxFfxg+HBe+9Hr6bobZixOXw+Ilxh5I1ey/2/y2usr+h1mM6AQqjoE7
k1Yd9UD6mFUJeQN+TSWRUDC4Q28KyoiaANGrc7DN1EfElpSMFUw6Ng==
//pragma protect end_key_block
//pragma protect digest_block
fr2vTe/1p7JlzU3yXI4qyDDx8vc=
//pragma protect end_digest_block
//pragma protect data_block
eYK1wg0MpCYdynwJCB9fOpZcCgPgkfjy3GTuh+djTrjYugkuTkW7DcqsheHOWXPi
5A1K2GlmRp3cIc5ff/ZTReOf3RQoevVsMuuTZGUEZf2Ev8xOvL8mgZRW/wPfO+jw
QcaF9+nveFObAOHuuJ4ymi+7nHtL03yKI50N0dHRED6PEqLoynP+qypoe4s/Ll8Z
LOFB07Qxy0tBJQ4JG5fSop4GSWKyz2cwGOrdj1dhyUCUHixLyzMS2uo4oaSkbLzY
Moviv8XAMR5L8RJkFu6NKrxG0AWkIXd0sHD/SKKZdLi/gLBZCgrWadkmdb/uTsv/
+5zJ+rXgRKK4mHdj7qRgnLrnBG2U+UZbL1ZKCXuQ1lXeyoYkDs/rH/Sr4bHQxZFn
hXfUXMVKSsv05wYHFhNaHX2Heg0jHqtpwqC7xYQ3LanqtoflIUbjWX/8BINcPqUz
8FAr9mHS2Hf/hyo7BTnzqrbWuieFlYduLCNJm7Kyn7KPegiobtMOANOBPiByJb5+
U7Fn1VZe2sky/DRueR84P2xH8FNHlXJ4QuA/Pray0MZ9Lp86ODu1zzzTHyGKH3Oz
KOlDELuuWIhSc8g48sYIEjbXbffr826dHQO2DB5trefI4VM2hG569ZCVP0QPHekU
z4hFHcUcKkVDP/LgViPmbqEVXZhUO0W/XT/mqY0tw/9FxOisdUoYH4+GNuG0Kzk9
1hk61KO6jnQpK0BXVCWCIJ6WcuW9fgZ9ca4sV0w3z7X7gWx81PS4KRM3y/WnIyTp
rhZ+dL9qfatJo4+8Pk1q0F7MPbAmokLLYJYC7PbGVcZJCV9daTc5jgaIIORS49nf
RTB+aktWo53DSPMCoX8oIW/Gw0FCvkZ5WtLNBlMh7pJR+d30rFO7x+p0BrCDrW39
e8zEGKheQ3PgZzRZc3Kq6rG5cci72vdciu2oNUxm+hnTAhP1u4CF4wTgcxfmpsGw
ubmZ+JT3FkyQkO/33NJkbHJIe3JJ1+tgdhfDpHzjDbaGt8ENQfBmQC5Gg9o4JDVc
XVK1CeugxPaoj6vtIHFyiXpcBwCXdLH/+lD9SgqyJwoWtD6K1l7L0bCrsDADFdqd
mOKZjB67/HTnMjb2lUy5HeBMwntjpGDsOxmQZNjtaPlb/sKuZoFeIDfYNbzQKAi5
66OQQehWkZ+vEbx7A567QsUCcFSSrNmMitgCS2o+JocGRdtanL8PcdnRDwuIGCXE
qlhl8Io0MaEM0bFWD9BIDnJ/+Na/ETnwHqJC4qEaMlIUCAsdCf3tfwBGbhscM27H
T+sgvIDLRM8A1QqMV4JCIuCBlznOU5us3jLpE3T19Zwxvn/geXQRYPB2KRqxYvwS
FgHO5wUhYp7oGTj7FVdd+6ITiDWKrqYYdA/ztP+mTdmU6nmmQJB3po9/bl/o4MNc
unxi9lDz5kMTgBJII2JNg4No3AeYOqg9fQB0gme/jM0LJ1kZVRQNxQ4WQ6j0MlHr
GEScp2XBJ9W4hRJTve1GqM+dMDEm9/v2MGt1FMVapwCkc8su1hduM97HB1fNfFgD
xZa9JvrGDBeOnQ6R1vzM6bh/rjCxFhJX1gc85bMS78uNmAcUrhm8PJfNxIpE6cy4
J2APZgkooCxSZJ5UZr5oF+TxhLnmIGdi5QG7uWPavCe1IgBrEcGqiQuXDlj5VJZw
1YjsO6CnKFb9/zuVMAktswN8erI3b2LVP1Jf0pCI5zV/uTKKUvrEBDlSqjardATw
FdXPEG8xtfFN5KcxQ6bNUvYs/tSHrqK+MhiVIJf4m5drYV5GEUl0O/ZsjdP4R2uU
AuO1TblJUjxvSRP7npxFVDeK2iH5RQBw/JU37A4tuFKySRxwF48bmdScR89Oh+Cx
tHmMIbn8jiyatAg04qw6T7XhUN6MSFvbfuQ2N2pJt3os0lMoIaYqmrWxK/3+ZBJs
l/vR2990a2soFwAMtwJ2bvKqLQ6DyEQXuqJjJIw6k0fG3mMqjOlTEvR20FkwZKAh
/vP7cC5IDxa/2j05F7+pZaWtk6LypGQv66PMmbx1Ayo+k3XlACW1G1U/IfxD6WEe
paPC4Ceh0CuW6GiOFawWo1srMFg6KTlpJeuUH7dO0Uvcn68F3YDiVKkW5cqIbm0q
W6h1tOOtD92npe2dMzMLyXn317OIA+bLCdiebpYHfFwScTHREUKoP0CZcGnMB69G
2j/LEF+gjlBp4UtsD7aV2CLjWepjL/SxspDvI8mrsQmKJUkrQSP5rMtmH5UyNP4Y
/iGjDiHQxJDyPXsZTRE8pWgLNXUESGOICwbSsd5uyc31bryVizA5uk6x8Dd3snDO
f4V1Bltxsgi4/384rxwscfV0qKen7W5LxsaSm/S2BB1+XlM0BI89ywgqjqI4w4mn
PuUhrOi4azCXZUJHTnmFx69GmPFpoHTJy+a6R2XI/enV6pWzxklLGxoOL5PrNGM5
Xv04ANITMnoJcVuzdLvhq8V6x9KpaEYgTJ18KPZZs7FAw/YMe4nvEqFfb/9uTvcX
vcKNhLxxL4AABohllvpZMZ7ERcnkEelqaRpQlcrxmt9LktecevvkuCeR62zzNsaD
Ya5dlXZEwFEQIGMNIVRYcK3N4jrOaeQNJ3RRNSZNidykfzkVm+XHNB7k79n0N5rL
AVqPk1zJM7aZjv2IcWe6rq24/6wmb2CqX+9EOZeMNavtG8TiyV8F43XCMl8KsMQg
E6nL3rgRVqFYnPXadrtWMXEYOTdDxEBu38/+nie+96KHcw0Efs048LdaFmVFaN7D
mISoYl8rxw/hiIKftaUYQxJ2pT1DrhnC9m2RCZp8+vnftDEYgMuNMizoOEzGjWoA
6i63KO9EdkmJr2ow5K3P0Tmaeqp0YunE0PfGQosM58vftwzcwxWb+wEYIjK8Y9Os
F/WOOX07tq5TMIqEmA0bHqXs0IecZ5gylJYqyEQM7kRo/uRSLUL3BWOQsH0BeTKv
edyYqhcgZL8UaroFd0KPyy8QQ6uj+uHLBh6BXJgnAQWODplxwVxc/TVTQfFkyeeT
KgfD1U9FShDrcR0flccKU6Z6xEnrkeU5A+2pUNGaHsiCg93ISadjylhF+9YSsTbf
FJZDyBItnvXFuqbOhjRTKzU5eIGU9D1oIu2RI9mRtMMPZ0Jky8kXeINNCrrlbAU1
8zLv8QNpuyQUtGRZ6I+VQegtnOMdovEdSK0AzKgEBOlmqg4fP4BfYXRjpYp0qwrO
/QTxnm44XJncPUsxMRcrxuFOsQNg2k482J7mOgnGI4BtLTMezd4L4dFndIgw/WLS
kHIGrw1dxBbnEEbHlEEnQqgRhSgKf7a4itlMQ/Jb7YZESmoW6tUWU5aZrfuLIOW6
3QYHAUOY/nNWfT1Mv7HtAGFbOP13Rxn/ovjspd5dF2+ytiWja7pwLWiRQbxdJk6b
h93ULwtMQG5C1SuY5LTOXFL2lKeNQl+UfcLpE3O91toXqahUFUwfpQv6KVvqZbm9
ZM4Sj8FwndLcfHABG3y2s7+P20AQnan7QpKbQato+w991PmC7My2ZLOhaYh/qC1i
y9lsfP4sFs1i9iGaWNoelUZzcTULe2l9W+4sU/BI6QFSn/jemNffdmwq/nBxofXm
VjUTYZpk+7C9493DbH4VUcPnATqDFUrogTVZk/81mDlBMzpjVJ97D6abhTTpmAyQ
SC4sAj/zxwKgtUKXP2VpRuLxEInoE05ho42Ork04KaN9RmAmjGRAY6Stw05pyCJf
0fnlMXD2vYFqDo3HeAbz46iQ/+yIZ9zN8lFWXGAQl2ZCJ0pMv6CZb/g53pDEnhqN
vE1IkfUKzG+gn6NMoRC+OB+HGXDevgUNdK7uEt3b33uh0ecc9bLlru0s7mye1EM6
F4YiX7ZfybqQRrOorPaIOQQeIyZ/Cvzr2fntc0EExlJiGN7P+lfmbppEsgkxdLL0
2h8RmRxB1nUAuEnKaSocZu1YWQyMjeTebpLxRB3cOEpvV0+L1fPxvUCpq8eQvPCl
o1jpFst88MAMKL4eEpV+9ugvgr/xmYvR5dMo4TK5NUYtKUbP4wx7L5UwR+u3aimO
L73hvlO+LMeA5NKhzX/zUZp4kJk0bR+LNn1iNMam5OO/t6GKVTQ+o0W15+Acwdwp
13fP6nubFBIA/pWd+T8ge5+MFPefbxneM8wbfwK8euxwxJ5DlrWsYJMH6ij/1AYc
1OY4A+d0d0w0RoMv41+Xtt+LlPgMLdjAgW8ATf0ZmWVfIc5biv30L5g6RJBe7IlS
2haKIWbt2toYQPZp+II0asvLC6xVx/e6hKDgrOGfz1oBB8vSxhYaeAI/GQAstChQ
SInjt/DEc0IlJ9VNmL6SzRmusNURvL58az2UEcD4OoxnDPHCAPap7NIGRDFuqON7
YJEU0XlKm5WSqfOvxgWjJpBOYSnynlYEg8IBda1bKd2x8E0NpqIvQQPvPABRSAJY
YOhHtCVapVtmp+rRDszvKBXFsUEv43hOB4U6xQYTddjl/HQKSpiqsjlJ4qwhFtot
9N+UUyfNzDX/4cwujJip7B9f+OTQyBIglRlZQAfH2NxZgA9j9gWmVyQug9HmfPVm
OSuKkuHepJLpVGOlgZRyD5zK2GFuWLcgxkQk8l09mHMZGjluitz9SZooEsaMDD7k
AvGF7qOd/E5EjmXHdGU5RR6QdZE3xOvq9ukbP90PQngVPGHIn6K4cwMTq9D/r29M
rvczAhXgLBvZZGBh1XJvhJFJoX6nmXhr6aSZIatKFpI25X3ZWetS0aFjJhcntJ7s
gK8vh2I/DM5Rh7wRZ+X0Fq9xIVn9Hg76NB3QFtplm9XYnpSv/BvRB1R9TTxrUHje
9zwWsmzbYqEPqtXZchLkGA/CCzq0yr1VyLFrmBOjDWxts88IUWMRH8O3YyNQNmve
PAI7m5VzOjjkU28/pcjC2deOuiK6q6XldKnOd5SePioWSRKlIZ8ZeOH0SIhicA6F
VyekVrJsOn6vB1ugLy7LOHhBlKgnixRxcTu2Qsmldp0L80eR/fjTROQtuiZhXcaW
CUNd/HEmoYkKBCxNo/53ZVwsZURQkUVBPmjMyfCPKw76r/3iCySHFiihWLJQxla2
LSMdXLiIh5V9IqELMbeSRmc2vMedOC/9BNriUUGklYkwFaWxLMCl1Bl+uDnMSLbB
XVBLghP7fqDa3nJsZ478o6RBZPhUGOdnLUdrtPAAQFhFmnNAHSSO20jnqds1twgX
pdYdSEEAMY4o57H/VLn8Z60n7SjI+4mjPIkqsW1CtJfxr6b2L6gJ7s7yQfnf8Qmz
8yInfC33gs/eTCP4g4LJXIj80OihzZBGq91WYI74NBwuAltQ2lRvtPqvWh7ScmEb
jWSydEKe+ISibPwQu8WVFka7I7Dv90tpMuppRR6OkEd3r6gSo9+sucVkCcaVu6OF
OtD3XCbiZFZnfoOPEPCgdOVl9suBoyOKLUcVKi74U2YJghLX3uMdefm9jn125RoP
l3OGYMkcVuljTvInRNMspDneb63c8eMi8yV+IYpwHbrWe1aTfERT2fkhw577dKcm
xVrssm7ID44lmTHAPU8Lgqp/nNpb1lETBnYgED2ayqOSAVctdD5j3KWWg2xKdmBP
+R1SzHMfFwl4442KiIzftPDYLCzGlgKSP/50pm1oeIXfRq4/oehjabfblJTQOR5/
Rhc/NbE1kYMwr0jmXJ7S4JDZqTGhCmcPygWkyDP8R10yTmj7JN9+hHJ/KcWUhCIU
zqVEoubHmFBOnOLFhzQ+cqXHB/yv9wmhNjexGZud3VpqvC1mLq5NBfWbfo6SLxD0
Fdqd1T91Sy1DeSYkmLxj0+yWfF8D3pmdMg/lBBB2PqGRn3uyfaTwAHGiEObDLgIA
y8xgTR8Prj7DxDrIj2szIYD0f7ph/OFwS94AZCWq1it8FuHoPbQzXv/kV8bJa1NB
W6V+N0qmWYHX25WQQzSrCapTwgfeR0jK2B4XFwjOWsHs/iakaoiYpc71IS0w3lN7
r5RtDg4aAgIvIw/pAqCViJYhEqso0W07pX6vVXsVK10puC1/WNo/zz47pwFFwa0Q
93RiG/oSpESW1ykhV3PnKMu44kNMCrILdmtzoQIDiBXyqmZNcGQgGGfkqbeYH8qC
2JvBjI+18S16OuwB96f2/lD9RtKrb0GLOxM8T+KznFIbMZa6ez6NJIYC2Ddjnb6G
Y7fKl9hcmvi9sjb2wYC/2wxTqpBgRX3VceVRYaOuByJS6i1J12+nayc0d9sM1FRh
pWhHF3JoeRZvSqVPQMdUKmjZyIZdr56eY0Kn9n0UwTHDyFwXnjsuyfaQjrv6TVqb
CAyQeEW8IfIM0Az3jcTzN3nx2kGwucc5tewMALb39fl9/IwLipiDwfJf2uELbZlL
5YIOoSdcyb59DaPDqnVoMgjokbapg2vub/Xs3aRpGNsU7MFD9TXbwpF9IZpzYCpR
q8X0Kg+BSSDgl2S/oCEVwDn7oYu2EMxNdKV6jhxcpG0Isyvsbs03x239liETVhLy
BnT+CGccYdp6Bk3Vfd9FipTWUSoNOE1z/xrX7riKrA6yVPMq0Lb6p0OWv312rKTU
JmScVVUG6dh8mlFzQEeIM7K7u8iCG38NvF7svIDXeIqWfdojoTzWmWRay/13DFVe
DKy8r+f7XVIv3eXD9fRr1nHdSOKdSbM0sgtOg/eCZsDkBXAkjeopwOa4+8i40nxh
8NGfzGR5sC3YZMUyQPtsZY70C+684ZRzqKIWtmkQPcy3/D2hGXOg6HDcjHg+CxJ3
/3bB12KpDcD3O9dxAtTvfF47rQAUjFIcqD/tBlnTzDalDmEf/Yh4kQaJzQLZQ6ic
8xqzSMp9JZx/XsdcJoLqcTEtIT47fwPY2ZJJm9KE2MB9CYeWEQtjlbkGaLfQzc2t
tCaSlVByf8QY9LsMc0gFzBBHeL1PrbGLmoLpvY7pc8b8mRaen0qBVZyFHlpMKfXa
8eFn+HPpxU2y4M9ULWpjq/7aH1cL0gfgm6ZDlfbeOQTMJraqhjyf+2uoja27o7uD
cR2X190jtsTjmFi1pdRREO07n9rXtODqC4mTMFlphO/hfGLy+LLapw68Hdyu7yzW
4f5IeBYhK9r6YFXOZfI4tZAAEJggUjWTjrgFyzVnluqHBmh90X/DIuXMIyjIsY41
pbxQx/mhnguFbmkdZiiuZJ/Net0foqL9CNRpHy8g9nqkmqslV56+4Alow9tbOAQE
1KdakiQ/d2iKepPJlfPOHXk0uWsi8oVQuPmw4uDzsTt3NThahzrQgneMYYLg3ZqR
qrB0S0m1QS0NsVHpHbDVZYMNS5cWeKIZPOW031MuZ7YwUHrwH3Rvy2Ed1ZJ4RvJZ
HP7cK8Oed0HHbvLkI0uuFrNiIXHtfNW/HDmbzfqKVlsuDi8epak7obYjsg8v38lO
oBixdSa2xCYTvLFwX+R1SeshtSuE4CJzhSX0r92cDHE/ltRfGMifA980OOIyMOX/
+r2cB3b6ohEmouXGNz9R17N5ou8KT4dkvi0XfE4C03Q/OlztRMMIBEpT4cKTSI4A
n35Ot3geVLyUXE5BSUHAbJogaqIe85Ikt2pnVvIQuFJoBeFhmchmv+PJMuh8uo3l
lXESlVIydhu3T4OUw8Yt0cVnkvlIOZpXx6aHBPeziU5bwfiLC7WXlz8C/wanOP4t
lZxeoztLexyvZFJCkUC5qWZOUrSdVDQosWwVHVJYsBg4s1A32A0f/VqryRUZ0cM5
FwfBK36C+HKmWSeixbpNvbi4f0VhfZ47gcEv897r8L7/+2Ve/Kl2vKtir//Ps4oo
3Fbzfhj+a64LqNpFTGg3TXp0DTLZCZJJtRIycJVjYXrTHXDkelgVqg5A+UGNJ2qD
tLWhRTsBD/d755A24KG+iKuWZ+GsL0wxvDBRsMzIEt925RYhULsA1SPLoDWcy6sP
Uo4JDv3wOHusrde51Of/QWt6PcHIg7oFUAc/56mArqxvhXFr4QaLGk6mIItrUYzb
dPdNBgWZ6M5zCRT6mBj/4GU3f5HGKatVy1D1ZIVDWCUJOQn6MEuoFguudKUYnE9W
GL1owJB0eOktCeLmS2DHknJgPUnctn/sIyoVpDaowskUirLizTMxNbee9aNPkZhU
qcGkgR7B04gZuDdvtFKFb/Sa+z5xTYtnQQ4ID7jtuoCHYOIH8LjIYf6gpBbPACih
vbTiOs8/JQX9oYXlYJYJzcj3mN/ur5fRai9xRh1CtNDD5fGsa2eyoMS6347w7plf
IMs3JwRxCgRyn4teiSQPUPbzysFYfBp/2P7W3IWeep7kBga2NdFv5VJXJX9Wx3rs
OdYntCPnj+aeK6WhoVQAPLHv0RbPoAPWVYWOjYy4Vnt5IO+KsUVMlRo4TRMm1fbb
ew70PjQ8TK0WTzbfXEASWXfSGL1rY1a7M2E8BxsH9aDqcNTMEedu52sVQtO1mEoZ
cz3qiiXeJmeAP1yXdekI9zEllNg5qJwN2g+O+j6Jq7EiiExugyUaoSE8eW9mCGC5
DnDeiKIEtS+8taLGPuibEbY2Jb8RKPsRX14sgxL7ogGpi5ZWjVBqqir4R8imVExa
2MTRP8OyUxz9cluBq6eMK+lzTNZ4MJqoI2WnOCt4shG1aw54c2FIpE5i3tJtaab0
Cl8tc3E8bc0jXKGrDdv2ZTxVcgALPW0MrGMqWJiqpsiyTPpGQvyB2Bk56nPW1J36
0grzgS9m8Q6WO3EIHGK/fCN3bJZEEMisxIEadm+ZoWCYNiJ6E46XLV+vSSPc0GG4
y7pNaOe/EQdgYgl7mH0zHaxsHVpu7tsFrRVksRsh8zvRnIdGX24JQRGyP5rAggdn
9i3w9BxNxGOxfi1W/ULY1qhsYJ7DGli8QcOWRavkPmFdYDWbMmueSje2ENkOLpey
7I1OnKEh3+IcMDeIS0G+2No6NogtlzGd1vnrkYpz7xcvJyl2gPYjLkaxycMowdp8
OzdViPE45rJpoQBCdKvjj2Rmp0yK+T3KvPlTeCS5PtutmIHAMgR80yO/Ha4/i70n
e+YTjirm1AMZO7SYG3YoS7szXf52hV1vF3+f7Hd0cYQ/BjW1N5KkgDJsJub6MUr6
sWJEZ7AHCiWLBEAff+WaCmHzdw/twOswHrpdXIFfNulu9IO9T1TKIlBM4DI/rMqc
6RyqQLWDXJSZyfWUnoSKji9IqTgixQQWawTUobRmTV5BJuRvXSeduLj2pT2zXz2R
W4ms8vJXk1MMnXZfyy9a3XW0aSPQ1jjx+yAocXtcMjAnauHQU6DQ/V7j/DDeIkSi
PdVpSZIXfC4Yl1RJRGbIaVlXFTwz5ASDlQFHLOROd28zqLt/LhfVJfsRnwwh0dXC
qHpXN1NixVkd+yJ4l50WG5y/4MiYiDNIfcj4zJ0qrJDMDVBfR39DyoHB1d0wH732
ArL5fsv5KTH55mkGD26dmlZBn/upLfAIiBC2txZDlOk/xpMgoLa289UM0vli+77S
y7x4jUXwrvGpQxEy9Ux+kmd7WEaWz8vl1bQCR9lDCwsi+IRd0W8rgYGac3g1IpVy
YATllShwY8n9ms8+sSSeeDoOYheuDA677ggK1cq+Z+eTtWtvGNEEbR1ce0Hp2L6p
VyS0XsDKeK6JZPmnNCb8Uz6R8TL8TG5Ar4VZfpVSmo28luqkc3McYFmEYu15J+8O
qNFQZMWat9K9y3sCUpM1lBrGeNyM29Sk6qxe+FCu9g9FU+vw4EdYlWdoC25hj9Bp
S1axtPk62LJufCR9z9eYlGK68dsy+4Pj3QaoDEK7xiVL2YeZOSnMzFm2X8+wqwSp
Ri//ujPlmK+xaTCL9cXwlqek5txnWBsnoEqsxmMRVU8Ig5Ak2TR6fRNBjBE+/J7F
6E1No9+e4CZcZYVw09VkF1+oqgyFR74OhnBL4+MRdybg+WF4UacvIP8MJaZSPUoV
VGIIE5eGO/eWvUw9LNnWh+oFficeBjlIHF817+O1b3aSbn1oZsrRMKWu1nDU5mhr
PLOb5x/XuMNBMHw5Jssk0r0CHhptYsxgJMSkL5JvDaeJwSyZoRI67Czfmcb4Wrkw
CrF5lMDKMBk13AqhgXX3f1WbRSPOjB5nEHdK9biBaMK4IxdOuNP1rduF9Z5acfEm
DV6QktV/RLpimZjcN3Op8A0YdLAeAIhQ7ezTYiheo6UoIBapD4Fio74USH/ix5WE
rT0v8Q8dUSEIC2UVzpHG/TXOV6qRdKpvJkYsNvz3U4tu/KVa5Hv0o4DjHx4/KcJF
TAtO/xyfbYsTrRoYf/Iw1Rb0pVWnYP23ZkqITXun43XEqg0nkecPi3MpCoJ4lSL8
JyA5X4+5/8A6RlwzS/uOMoAb7zmO/WOsHTyFAZWxLRGtS/3kCDYQyoPLElkCrXec
KlhkQggM4gadxoru6tQDPDDA7N/WxJXYTdz+juLYttl7yZ/4MHxumhOviqR4H5l4
IzBVbl0I4E7T1u+fH6gb8CZ78960VqspjU9uYNYb94fe1CVlaJcxFBgmOHOmyEfj
kc21l1ega2+Sm0rqdQ0nPkVob20ixPqB2c/AyXARPJ9zgYQ/cRPnlBleIyGxtksz
QF8J9Tf/h02N/eBMhZxyFDYTZjlhiPjNrVc1BOxQ9BEV5XtewQlW2mn36PqGbQiR
GsJJyiVZX9bBYfJQ9Nis3jfc+6f5G7b9YUJ3c+FrxIz3PaGYnYnKyQMOjqUr6Axe
ogKCxwdPieQhp4pNM8oUwFLowfkSSQAx8GZdB1oF2VO07zFNEnVQ41RWwHb4fzsA
drKe2oDn7gm6py+GngmsE79aOaK5jTqxN0jfXD86gKfbJZ6+ClbWU1OZZdnw1ERI
we8w2oJODiYlHQRGwc89OE6VHM+28UB/bkYYn1d87G9K5qmT/Tx6s7040xlH8UGh
Mivv21OAaEs/ANp8G+K+mXdZZJAoemuEq5ZkKlBgsx2pJVtpvIcwMzif+vNgjdD/
3jUMMW+K0i9cUil/2qyTa3ZF0w8HlWeYj4byO4LLbTnYb39P7FwEi2XVupzvSS1y
/KGOEKNLdarerE4TsL2JXnj6MKojQ1Nlkqi8Uxiw2VS8XHvOC1bSd+iMFc3QNZJT
nl9Egew0lETiqjOicPJ75WG3Yg7Fe9Ksv+mXpHPc8UFTNAHOY7ds/uGweXw9I8RA
8+K2Zl2o2SFdLR0jVDe/sKtc8lwW0nAf9W2GXd+Yy2xp0U8fvvpXCVJdZtONbF12
mO7/5q3VNBqw/MNrMhPXl584tHJBBrjQGiriXEXQEWGh/OprdLVnlrgJUZFurNoQ
UC9QtXSVmmwCGBP6F5GDm4rpg/iuIb+4t6HnK2V6sqFDWn3oCvcySp7EL8UfmQih
lmEbT1Tqcgs27lxziDY3dsBwfqAYXjMEL9+Rq4iYy9kywJAJhXJqwAIZjJgx/Up/
D47pVx2ZrlUTTCPcmHONYTioqoCLYHilefawaLXzagYZXACSC6ZBI/cYGMsgyuj7
mMJ8esmYvNoG7Er5qjNhFLE1sCfmHZYlvck2R/77G0m5+8hzRvsQ98g8zGkW+RHe
87UpUe/x0qxV3K/bnjeHnDM5W3ofWGNbAJAvjGQss2M+FIIBYKtJuh81hXqa6b6/
yd7lDBmiF16g6Tb+7j2p4unDPAn/N1KNUIbB++Jbk+Y3YwpbHK0mL2jGXeTT5pmP
3QnVUr6dWMMNrpm8D5+vD7tsJq05YOPXAaDj7xLvY7vaxdRKJei6wotIHR/HG6JC
J/5iv1pnEcvVkFrnIVsed8atoltc4YMrddIL1DcEeDdS83I22tn5tAceYy2b6d4W
Y7cfRY6wYCbIzWAa47JbsVX8QbEFtTKBfi9mUjE57cbwDk9R1CaPt+SimBbUXP9c
quMzdxfpVYNKYz8B+vgv+w1VpxnF+6zPaKFUeTn39/SjcBfq27LQMyhZChX15o8O
f+gg8e/6AYgBPqdbg/UAiTf4yxjly1g0i4CPhKl3BGzu3jxn8j9Cb9mN1W2u9rZV
EDo/DMtzOQr66d7mvgjgpcEcoTqNaLqpTo4jKuw5u7EcVmN+gr+XghzSN2LNSZeP
JHje3SGs2BLdg+4V0GZoqJ3j/ZtrNbkk4ZvsZu9wZK1Fgy4kw17q7pADS+mMamDN
msMkzZmizI1Xr+QmDDWM4NV6gB+b6IxkkyGayfhGuuL57Yo8I6iLSgYP/tPF4mTI
GG+JoQYikZMo1Vl8INCkLES4Zc2+My+DfwCqKZ3HQv8ZmZG8Fkx218mpOGFKRMLe
pNBysb3RNVI3TPbi357rhgdg3GrjMCCAIySF7Ku+r8U2w1kjVE3cxkbPbjIM1+d9
RjSnXcL5N45ftE1QsHEZPd2gT/R0nUy10aPUuKmzfcpYr+8OjOwjm9ElPuiiWE3k
eOSZnFwHeuglGpCaJzMeA2HEkp8OUnJP/xv0gfHLKggrzonXxveciOoUIhDIyrhR
jH0SHP3zNqk1JVba+zWE8stEeC5Ye7AMoHmtWxeWVHKiHyx4Hez6sBhrVf/KF8Ub
QPL8ix/L9qs5T/qUzXHp/3LciZmgXHkRYIKgVU6H999FJm0B94nqzNr6EsTj1Azt
+ox/nruhm88LlzoRpl6bzS3x0+f1XTp23hz1wvh96p3mD4JxaYc8fqFP64s8U9WO
d1QF2/eeiylAQcIAlavDbrb6b/LhtJgfVMcacfGvDafE0foFUwAOOZeynpdbar60
0dzuqnk7c0AgmbkdRJOWijcG3b6nWfkcpEEWqu4PqXk0Rv+LqygeX+P4pW3N0aTy
JY0hvVM04izrh0lAjZNodM9q/d4iEtLS83bUW5eB8H5W4wSO7UkdDy85kQ78lGdD
TrRiW0P0CJ/n1CnyZ/BLb/KHUNS0T9pKzG7WPv35LULDW9O3bWGk1qXuurh3Tc2U
25K9NQ+5oDk2GhONMRwzlyphQ/p1My5AkHtV6Uo9FbjejRq7vq0cQI8c505RSXDL
XkBQn8cho11bHLxLgYyKZDuu/fOvcqOvviB35Dc9lLhXu6cSxvvEwCBvVcHMj+1f
uwkWOGWXZMA6hRYaZkLlgdlYQ/tJ1CVIfQGtizQ7G7xx8N8c0E6msiFzRRI7lRPO
15As/ZDXq+Qek4GYP6w+vZlHVkHMuhx23Ng6HYsoAbJCmRoShskjTrTBuFWgHiEy
n6c8T8bKD9/pI13s/qC1HUWs1TITXkYa/ctJfa55TgAN9eNGz9X4avyg7WEckcrO
+khcEfdUYvugqeHyZrPAYDSzpgyb30FUFNaPrt+ahv4MQRpdjSUT5r71aRwIu+Ss
U+H34oYzjAECZGNTSgULaBUtgqdyN3YbhJaeCB1EksBR1V6yt6WrrzSeXu84d/8X
OpwE2WzDRjdtrpFj4p0Sl2dL1aOPc01wJkOOYtBsVP7MCHVbNB97ZmDQzh99Rj03
MzqWloDK96p8dk/xRX/GeXoB4JFALrdd8Ud+qq33+srwPSouqACfwQnsCvHbQMZr
TPsJ4F6YAsP4LC/LgXdvy1QV6eKJ+a2tYO6zRUGgdm8wD0g1kmKVc/vTbAeSQfcv
hQT8F64Y7KV38khp/3YbZLdU3k/PA0VldNGOFTOFbyp9wB6FXKNaLLwovJ/iGsrm
GvxtdHSV+jG9OZeHLqhp6UnGZQls+VP9ApglS4GgZm2joYtJ9r2Y0l/uLBv5YryX
ZRXNhtPOTlC6qldf5JuY31q7F+coG4LENo6vHjU0SOwYtXwFnUKdVmU8+H1D3rhr
wSMoapr11e5S/516rD/ItNk67Zjlwo14TZAOlFoHE+dtY+6n4iQueLgIR7nrWwEj
N5F7eAtefXLlJLEkXlSnq0fBZyd1h+hU/x8KjimZap2l70r9iYzRnBhl/R9Fse2t
vAwjuTvodgSChly4nDXR3rDTN7pMwGwIuaPEGX8O6t28P5tNZfgXQFGGsXTmTVKY
i2OQf7WbaM+WVmjmZ5aFi0VvhpBmncabKEMZkbknH25ij9pkzQuLkfzvKToo8Y3L
4cdkHl5PtdgMv3mU3z71hw1Fvc3MMLRWzqtC9EQB9aV019Xh84UsyYQOKNVhsHmK
L23w/8T+r6tlTUM5R207lw3k/eyQ/cqtqq9bin9cr0w5x98n9M7zoa37BFeZCDnv
ZB3ueXzfEBhqmjDC0yWaegwofnJ/bRDcp1aLeUZ+B61H/tZrSWpQVO2C9VAS/qfd
GHux40Ch99RvV6H0wPo8lZEFtiAPZ8vk+LY3SwE3LaryMnxf1X/BzWNu3NyHD93+
XsR+a0DkAM57tWLw9Uw8ah9N+x+xv5UY3dWO3bkOinamCQaV551LW7do49GbpJv5
WjT/QoH98+7vMkBiapNecnayuLXSfLXbStS8Y3kUWotjQt/ZYq7DnTyKBwTesnJX
mrbWQ/yFu76yEKZ/Jr/IwLBpVoOGSyAQqeGqsKUUpsYUGdUVhU+mENq99TS/rbIK
1KQwGWZy1Eudb8uoojy+48zsqkYZd/gW4a6PgN7HerNOjO3aeRwsHYR//qfGTByl
cJBwWjrxo8Tw9kfiX9OVrxCoBLscV7pQoG/n7GDykbMhkoEJCUKbnYXPYA5JmtoX
Shxy/z2v+V2rnmwscCNPti5jm9Q9YYrYbGnyP9i+51oFJPwR6i5JvR6mOoe+uqgu
i3EaiqXpfUZ6QSSaLulkqOHjJUP7EdLD7FsN0DlgRnMaFE93ZdLA26g/6rFbzQrP
asIaZTlkxmvhrI/zm9ATyiUxzP+aNXY93QBtbo5sTWcwuFEw/1kXCQWCihrzbrvO
Kz1C76GecJsaKjd2HuVMSpE8H7P+R6f7+nvIJPNT5WBw9hPabDbWHMfvw6w/IfYO
/OYA1CZNHgTuWIADUwnxd2md11mwE5mIwPh0rn3byYVvVaaL2TL7vSNfBDcMGLjI
/NaSaFn0+MtSDjvSUJBo5VmLBRmubyDQk5odjfCyL772+qj+sH8081s15IvmdZDD
QRkNGpF3YsAhoYz4/YO1hpvalYuFhOXKOe7nVS8be4gTsg2LCMpOn3MZodXjFa3z
4L0O5kXmUSmp0wEh55Lqdlrjp+NQneWxzKlMmKSXNLSrh6X7pNjhk4aJVqtV0MrI
mZGaVoSaWkTIAjwNnNWNgdS+O0JsLFecmI/on9ytDnVW0WFPXqiBTzqpdduh/sqg
3J8+I/j2nXCclYXpyoRpIQpKsJyc698M1Q8qAxVZXHGLPOZjRp85z6HUAOKWeL8V
AIWhNUicwOLp02QgHTvKMYJviUpZH2OAZALO8j1EAUAnDymyvr/BT2jdDVdcanTv
98yUpsbEieNhhYr3kLnwBUCW6DLKUITdrEeVcCTjzAgdq7Xxu5OBmy0yni7yTQlM
ef9o0Tjn+azzOKCcPHNpRPJo6PrIIdvnAiGxgntU4jnnBjdq61iWNMqbqtQibvBf
hKij/QLekePu5vvcqLBeLdL7/ylRe/7W/yZuUMVLfbskEKlri3kmv0YePnhlrKTV
Sj7/E7QAj305c916f/VHGDC1bSPEE2nvT4VDM6URfwlB751Ek78Nh8XJ2yoEGI2Z
H2CvxvL8YjKlmuvmc9O6EH9ubE/Opka5Q2OB49DDTW4ap42hltL3GldAOk/BA80d
eeBZbqZF2gO1Z9U4xFRAu69ir9srLkRzAJuHXbtBYjxzDVY51gn1MCiH9a3WuJQO
HgtSG62U4y6qoIoh/IFlLFg5z4it1rk4GiRnBC5D0ox7Hc79OKRzcrfky2EZA5qX
e3MwTPCzY6r6DpWMgZmOgK6yiftLQzKcc6+g2Nfv2M4BCDn4hbZbmlFj9EJDuj3v
+djsXJg+I5y+U+AJqebFPCQsFQVeAc3EU90vpbtTW3g88Ya7yFEZipXz/bphSjx2
GkpImfL7yfBV1kWv0LhzQXNNuttXHyJhO7K5OcU6yDZpe642FDK3dnt+3+EwGY7m
tb07QVXk+CnCvWTyLZxqbLkdQAolIddQybC61biwnt1+PjIO6aDQv/IVtKUzw+T5
ZY94Qi4uPw5959HYuP7CoWgmAkeO1SWhZCljRZP58Yt5nf2qLvTanYKdX0vHP7Uv
1o4xFbjrfcygfdEnO6Jd/e7cjzklhUwe7tWrBiONecFB/py+2Ip+a+/KJP0X+98Z
SxolxruYzNOtRzG1XtJ3YM0jBA7hRtFtly9Jv1nAcbU5Dk8WL6+SvcybISMl5B05
6ASW/pe1zG0o3wuF0P4lpq23odvddZILHkwbVmQ/vbMbfdcXpYPU89FdpNZ6pF+0
lxRyHWN1SuuSW6ybvRs53buwEbJ/mu+j3SwZrIPltIgT2LFEvzmSYpc7IiOBAZNJ
4gRS7Veotp30KUsBKMltpewYHVynYdQrnkS9Cp/LvbyxqvDIuuZfiRmTJicdeGKG
L+bsvBXIlhVjBjMeF6u4MShpaUY/HiS8s0vwWOII5WrKArTJOBcc4WPg9entXL9B
qc2yAR9rXjK1Km73fwwUYpI3kdTAQ3aGSMs0Uk5VZ6F2Pvf3omzA+8dixkc1MB6w
LoQUfDbElTYT+mctUAUrPQAtDKWln6f6hSWA6bkXIFj+4kK1A8IccT0Su3740YEE
eT2PWI7GlHJoKUJvm9acMoEidKjHbE3uvwU5QexITPwT3bJUT/yQnipG6qH6Oi3O
DWpHH3eWUonBR6saXefqF6qP36phQ0wryAJEgkeLNr3G5GJV5BrCY+/n67AwJuqd
S3W+rXLIYpz8Mxukq5mUcQQcsb7Oyo+gMEHrhtoDCrrooUQfqLaSLYeB9rKuhWTL
vmILzSMjAJNz2m+D6P6P22AEZfel8NNsK0GNYgT0quNzymoQCg/cbSdziVcNtLeg
TL3X7cwRUVznIEpbub9EaKDLUmqUYYHkZ3NWWa3RrF7J8FVi46jXVAkYeAn63dpP
K+lyvhkjNY72cqOXy9FRgkAF4HYB9KnKa0qZnOP03s5t7e5lsSDYdsCA07ieVxDl
TdKOWxZqPFK6hOWdIz1/LP5VMz1UMm1YGZxzRTQ98E78kIkKQSiWOIMmqC8o6Tqo
wv/5joq4NgNcdKaQXZFLzfhlWsJYFk2PS8i/fV8FsPOt1k4yw5J2eYqg9bs5r43J
G1CtkDcWQKcMxTJhh8ilLq3//C0nFdNT8EuyvD7ox2dsWcipcL12diPVMSih45Ex
ufslpm6ADSZca0x+OuX21BlDGixxBanyXWRbgOZzNejDi2o0N4jt76vwNVskKSsi
dZO8ZiYMaVyRg1ZNzwg8hl+3Vk+B6kMr7mQMsex8phth8aS8c3RuOoPrBvioR5Dt
8fRrI9CWGPrO00ju4/qDqATPdY73+tv0PIZovZxZEsakkRiUch7ffti7fchA3Yug
ME8DNd8mXsscSTUYJ0TWzYRrSGTMBIc3QtM4djd9TgabucZ6irvNV5ZD8o7/ZhqT
P8ZI8g72/Iwjew0yncL0j1V/swzvEbnMJgLVWspnVsAMsbdaLdbmkvkoi1xboIcs
Thp2qfrh3VDSQPxa/rwZ1/jJH3ZOlL1UdX4EcWV41ykp2NKuFYoYw0qKhZ609BOh
ulciMbFQPzYMRbqFXW81jkH0bTRVqaJDHGI6O8DHmVlm+xL44v0FaTNxdim4TxwJ
FO0KCufD+93hhhWp/uFgTqjpY4LAqJ1aJ/KSsHSWXQaRUYiDFDm57NpzdNWRxTd9
MEHp4gfWtE7J9k0mOk2dLe6KYD6v3rWWT1NeoO0wRGJdOf6glxDq/+NJplXM1o3k
lN+gHBi8VAS6Q9IUK5uEIpUmyVlkUaupqEnXKNg5yBPt0K5I+ECWxKkfeURQ7oAt
CNBkLBj6WM3eHRXKHZ6oNudPLEx8eoStIL0hZcU95cIYCkaY61hFbRDfGAt0GkIw
InwlmUBbrI4LTUr4lWoLN0sA8BLUGD5ZIH8MmC2EeK5TEp9PCXXBiPq7wT79Ay3a
cAZ3gqtZqDbAReincgrYxhf87UyrCe4HGvomwAkGDIS162MNRJr1QDlOaO5egaHC
6PggbJrBqNuRfUc5k794+VqfE1YcB6fjSZKMGnKwhycRWt03NnKLgMW++QHMDn0g
mu++lAKdat5iyRpKpv6VZJSG8jkxWFFtl8bckjaLyAvUigmRT0qhIvHoj7pTF1yA
h4ftfvM4SV6OjpMaFC2bPtLf6l6hoY3mEFdvwHQZ+bTRSEmeEpm0tXY7E8pRWu1M
29KkDn862oeMp99Ic2PlZdTr8okJELwAwNdU/i5IaAiuNWmRJyaEmF34fXFsOVvG
8XbjYa7Yl4GU9jhRZ5VolDwaQl/8bdrvRXB542imYye0dUCsME4IkGrs4zwMFKIH
ak2/x/FDuH8/GeIuDvmbXsRcawoPpPTj697kKlrUTLNg+2c9C4mxlyqG85FM897u
cqnasp+8W43t5RjRLbF/fiNzWsTmOXnoZsHUyecI7uZPSK3BfIAhhvE+6jjNvTCu
aJjLLKvExmog8Am+jPrgYVwpsBzgSOIrUMyoCA9zdS3KW6Uht81QXa+gqGv2h0TZ
WHMrDgobL6HN7gNoy4G/aJVjFbxdLk8RyiPC0hc22IDyDJutvatPu5VVkzq7SIlq
hzJ8IV/AXFZLUEDRLRMjyrpmDSsjdyOPSwle0fB+mQqD5FQyZASFt/PLUiVvYtuS
r2MAXGV2eQc8TRgBomordLKrXOTdE8RVB5rbXGXe+8WG3+MSE7xN7a9JFQ73Je16
cvfXTQQNSHeQLh94i8VIF0vJg0mbnSt5ZlPC17XyeXrdoHd/J0wvaB5XCNNkj7Gj
kwSdMFMRBex/ANsE9cG3h2Pg7UE/FS7DCLKX8pbx1TZV2f9V6q3LvP/V38Y2S3r/
z2QtruCQp1zXfATwAvs3v5BmhwsiPFlYU5fkaB4armNDkjS9NdBIvmnOEr6ZsnoI
03iNGHT4/g9ve3WsrXg/iAy0K07GPQRPUnZsDCVqkwp9dvjz86Xowl4y2kR1IOq1
Klk7bPCLeQz/OLyLSHv6ceAUJxcqLsLmaJVOtUx516NUkl8gUMDCeBjeOMmJT3jU
mi7sQiZrCOz/tMu4YugWzYeLWXRkQJLiR1YYl2mvc0k1BAur5yRfd+XXVJm26z0B
vRN5OJznjIPsN/b20T7UBBroOY+D/kLGQC1B6Uj0zS94m0m4ALnLLa82LtAzjRmC
1ZbSiOpNknWxr+eymIsl5eAqE/s18aVVmuGvYLQg9mRK5tafRoZLVJC/+aiT3cF1
Cm97oYrYTgq67tAmbtYQpFye9W8gMkgyu62CiM4+roQnJd4rqRF4wqkOcclOSTvL
sIKljn+GSwLSIVe/0qjO0i87WGA2J2C6dyh2mmS6kS+7yNma7eSqGvZ45GQxGy+m
gLZEFCMDiHWzcLwk//mI5U12RcGQda9WbL+r+XP1VE08mAkuj7UzJ6LJSQjpKmd/
XJC2/9V1X3LJod5ltM99p44jZzjIXzzpSD+AB0FFINc4gL82o9O5FLkYBu9FxfUF
w8w4GqhqzNuAyL5JvAB/V7hAT388mPLABDmTDQX26Rc+iUCt7PUhfstxh07LjBMh
jCb0PSMn9gX1VlqI6iAl+ULV+z4kjeXv3IxAc5vMUJ9o1i6aVax+Rg2uiRBkm37U
uMobxAf7+4oR+oaHfF13dzAlGbv1i/PBxOOB/RoK5Z+9L+MVwqH2dP7bES79D80f
Wj4GX/pf9dv9QnVu+69m2/o+f3fmDrzWgWr5QtpGm79bg5VzlKXQJ0a5OWfmmyF6
QCkKOi+dKWooO7wBU5hIBTs5kak1fZY7WodMIeVITFLNwm2bbY/dxi83xgIeLPmj
XZb5MNP9XBFNepXC7+xuT60QJQq31HrfoiG5Wcls1KZnj+UcCyf0yPnEfZvr1AJz
pmh+nxjB2YhLw631TkXfRgXpmsyvA6XqzSZd42sfBAe+pxS2VynylHVsqo4vyfL0
F4CEA4g8dxDczHBw+ZS1qElUoGt8blaJ7qVjszh6w49VjEaze7CmZhITO0njCLBz
CHuOd6hls76sMSbhM/fmqaLAEOIyH0VF80HSflNLNIlllfntXlen/WYY87pUaZam
ORfj/H2lPNgQDgU8rXjUDVAumPuRG4Qsj4J9ZIQVISFjaPLIkvNa7xCFqkcw50YR
0Ns/T36gncXHoBacdxGv0GTz0OmMxeCF+6r5UwE0RbGYSd7AGSmlFnQl8/KGyNDG
Njetc6HkgVYNmDYj1PdRfYqKJ56zq/wYhd9nklPwuioiHB5+00XpknHGyytOTuKG
mHdttb7KId0Wk3rqPO18yfoir1gHxoNrQ3sZ4Ep8LDqra6Dg4C2GooS1UmwGh0kA
AwD2pKliC9g6auhuy6ov0XCedAdExA/i4jblksKrvSheiu3lDOQ/mx4CulWF0R5j
LvBVk1EkqN81XUW50pJwmN0rkiq1ROyDB9SxEdfLE7hQ3S9uk6GZ8+2IJQHNNQSc
0GwiF8BjqlCQWfTwz7zzjJGXXDe2P62rJxvviZrS05ifsPEL+YwHr18df9Sq74Rf
H+BhY8+KAb4SO0TZJQlS/r9whSyS2MZy0O94aW+BIift3Ah793fZYblfjuEj93m6
4B7O7RFvLKtvvovEQ9ft/8Jrjkoj9ynfUsLWFot3XaEbJEpWjEuWl7mL5NWOIl8L
emnRi1AYyiIPDcBXl6Xi7wWYOCz/t6VC0BBx4qAfKYkkWCQUhNvMhs80E0w8LQGG
EzFz+O0meWt/xSI6wGMmdbknOD7Bokby4KBomRoyWjbmwuYcQcrSvePVs40n8wjR
iiRljsHDIEbmSm83SP6CD5/eRwajDc+TZTzpRXwjblCaEnQokUMo0TbW0VGka/SO
fH3kU66gC1uLpJmfxH7sUQjgwZ2e91nrQedH2y4Z/uw6MtALBst2jWWSX3Aosh+8
ygObrrZn/vwGw7EOaJdU5JvZgkXZ9O5xaExLGNS506YcvrwIjtHqh8q3RATxZIsC
DeGyKceGdqfWdPxM3Px3slO6hcb7fwgwApPXjW+RLuzgQOQXs9DzYyekJvFVR67P
dwfQXZ/c3WHWJC55K2NFDGbjMKjSyUul7XjPhpRX/7OMeTcnooe1+Ec7o0q3eRgU
wI3W07GCX5EhxSC0ohPV6+x94zG7qOEUSuSDfupBhhttAcMzUAS0dmIJT8Tjzev2
WxD5i1JFVTbuPiVnnwgfU+YxI4gr8W4dPp7y0+YgNVVzhuANecaxoMAxIKsG3zGM
zNkyCMGOcyev8ioDqFQcdpjb+nmIeHSHi9byMWzS0ZjHOvb3Y/lx3cTCAiPVIKG/
1IwobMEPkh2WUAXjV/2ybJpL7nZxNjGcBzoJ6EtxQ4s9iBagyR2L0tJSIuHjlI3q
pLqTHAJVpFJMVDkNB7iJweUSvBz+KjY/D98ux9Ti+0Q8URE3sEfYyZ0hkCkEvvrk
ykcHTRGdtoF7ajitxmGFyhbLevSBMUXHe0SzpctbCpF0f8J/SlJVG6OISXHvS7V2
YpqGfXgkRwwKrIJBjkQEAar0FEEvtXewSCkm4XsTyvHgTb5oLAnM7VNDBoTsOLQC
r7sI3bD/cY5wFSqhVaOmeoeypuGgmz8eyaOwHkzHW6+cOEAAR27KLsDJGdY6dH1N
ntBKnH2xZiiJrKHRs94HCvK5NRlSaNTUBuysKwfiHKU6ywFc7iJh/8ecBy/MXvOJ
w88bAaH1jVE0Xr2BxRuhr6+GBWHI/HqJuGiLjyh0seShvR/nZyDMkdN45Ym7RYL8
AOiMqk1vqZNL2sNk1X/HoIUvEHdRB4WbOyGM+ooYjcUQ5PTrxpup6zUH4vWNLUaZ
/SUBO8iXu3d56QySpCJlr2ec5Yq9iGsLQV11iuNDd7889fEuQ3hV0W3XpKSYd5Lf
ViDeoYwERlsRHaJl+OOS+uH4xTJCVh+tSXD+32hYjldcT4cZxD2FFNM1mxdVJnbr
JfgieAKvfcglkJFd7Z+nQhBCXOwt3W958W7lNMMzOg+SoaIGQ1KV+z18ffxXDW3r
01WnEUxl7oJ0XNyURwnUyABUg5Tb06Ey9JPs2IrDU+TqKkIj0O78yA9iba8HEV8a
YJ/3uZ6j2zsea0yA8RvgdWDeUH2m3p9IPqGvko5doVwbeYtQhuVkFYkiXncmLrsU
UY6X7iDn3eeP2aad68mm+GZqOD519T2mtAXoSRSN7pVFWZO3VEUkjwuCCVprBDRM
OPDBVsLhni+OgXRJ8OQop8fUdtfo9IjwhAgkEteclYo0ay+MbqyU0mofGfSbxISN
dA2jOBu6dgT/4HDDk90DuX5TM46NMtU7ldwLyRBnK4gia2pbeb4iAlSOfDStsWJU
aBEsYucMXRtJciIiX3Ito4UHSrv0KibRjhbSfNkTTsGkSjvQKQmRbKT0lWjv1KUr
9XbgIcOC5JrrvMhntKi9iFv6tthCNglWLAbE4mLUFKy/HgRJyH8NUL9I+ac22KEv
sHlaaTIkTQsC+audELorb2zIrtlha+gT5gWsbXbRJAJTrChgXPtH+x1SX3+QA4MR
89wmF4quRZVeAAjWPNr8Z0r3VmmTGcWB2blADxRRPYw5CiPZOStDYiwrFLNZ+pIW
Qx4K2U9eoHIHE8uCbmts7dRkQX3z4KGjIkVmhe6ifN6Zufp7ivHNoRov1RMe7Syj
s5xO+JAHlkQxDjmLPsr3LvcpGcSCdBpeXKwLjLCH5NIzbyfC48rge0RspR/hxlwt
nMf1Lh3dZyujiIhabyQzWbjAEt1vFgWQwHlty4cAXnKQV7CujWjv31wrzUX15MNa
wmRRUPIF4xW+I7ysWDJX68B5c4a0exekY4FJ9Pyo7duE0oOyVSU3EgBfcOZu+AJI
k4VwFLeJL+6OYVVRGyzN5vwfIgC5mmLzTL8jqZdgLBy3tgncgT8axXMc+93CDzIT
EkNjmqL/LkVdTKz1OyKS0gzgpiAkD5l09Nyb5OC2Jex75j5KBtTDGog8yJvWcYIu
pY0VdxBPBeRV9ydVcEKlWl+LXwE9cE95IXwqzOTyb7Ap9g9oeIynDXiIycHgNZRS
0OERJ47gSzmmFl5FLzqWCYW84M/21CjymshS1nUwypmtibdLFck50y8orMfMltEK
0yQ3ota/yKZgkXK01K9K5JwaH6VISShg0daUojYk/dmiS1/E1/XCr0HFrJkZgeYu
opwm4QDAmpLpS7VT2wvBldsKfnc0uH1WeG9t4zOXY6Vl52NKezrd9RD3axrMuos5
v4zfkMUjCO69JUMHq0z6dZoSPzdVSR82hvQzJPoYw2HrNz4LTBbuMtZThOYXXjmN
YaItp8xeilrkaDfBPnhluRvwHEAHsK0kSe++onJUtM5jVABZxnkXpDNyzjeHetxm
hYg3SpmhwHXnZAO+hCoQY8WVhjWip/QA8umh0PTC+aUxFknxvabxW64HQbi+CkEC
9QkJ2aYmmJckK9k/7zO1pd9tHgQIxnLo6wEHAWTTSi5iZxk43QVSgKXWqQkP6eI4
rfrUGDK9zcQyfibwi+DW48vaz60NPF2g9TEcoEDt+0zHVeV8w8stRqOF4w2+tkud
OCOth34Ou25jLFGzuZmhrP+0pDdjLFLy7JjG4nF5qX6ePSquekJRsu2NZVqbw0Qc
5VNyOurWKcVBl1R2UZFjToCRk1zndVOkIlpGzIt+KRIspw4BZ9fLmc9u2eSFkOoX
rRdFJMDRc2ed2nvegeUTSLrAKucFb8N/4RLlbomMuu5e2H0EMel7kt8Z/Rz+v4z8
6HPajZYqUdi7p/EjMMvEIery3rBZ9Rhx6sdM1nDlGx25QZ91P/DzyD1fuW/GZuf3
9b3Vk3OsUCA5J263cYl7ilOhQxwZykDwmTl3YxwBRKm65KKH8sj5KMIJ/JLkGkqs
sTZM2zvuLagJxVTNO3tTINXu3om4g2xDtUydt/9ysvXBniv9eu6cWl9pr1BmgBcK
5X+n3lhpE5tB7uk/SFiBpodAQgxuwogZ6dx3RyzNA9LVYE3+AI4D7zDT7dofwZKH
sCm3pkC2+SdXQpaExZHwu+NQO73iMaClbIidThy51PMJi56pBQFSY5OInDnLwrMq
nf0sXvdxGHlPaG3ZIJ7XOGi2lHmfG01toEJvq6jlJPGDsPCbVduYvoqdMXsg2gMU
lU1tfIiE2xrkOvvkzN/OC6sC5NZqRbkRku8HC7WyEBmdnQkS3J0RGrOS25dhtgtF
kM/Pg/Jg56xgykj6bvSTE1boTdIJXpm7f+V57YCR5yWj74adZ6Cm7hMWdg2k/ieq
X+dVk7t6EY3eHkoNVCGP0nQsPGF/0qr+jd5TEoC+tNOEUGgQcy33cVSih2/cgEr6
6k0SoLv6UZbNavUeZliKzNdlIYjWciAAzIekb/b8V4jiThXOJAcGbLszZ7jsClAD
atteVCTM42d+5vb7uAjAIa4eZHvv5wvy1JHxksUu/QIpHRV5P4/9FvRrZU5OlL8Y
C1bN6MhTwqDdAuu30bIcvM6ivmivufXNq4ruRYSZ38BHdeuzeFHDoMxcHcZ+/k08
n/z0Mf58xww6vU1Cik79yRq81iSsYAKeEDbPn1PgrktfrPkA8o1th1xyn6tXrvns
rjpREY6u7rpGE02nQ/CRqU8vwOxSMveVTuK57pBIIAW+iGG1BUNhTBJr51FpZICR
qRkvgCmZkaIekRt/5zHh1SYIBJW9aax4ZicRM3Bs9hOC0I2eGBvmTjwis6RC3NJl
3+lDdsG7QwR+yJ1gYAtgyXmU7LCouCNKTrDBdDaP1LeJdhJ+0JeXV9P/UkwxVNpj
VooEeO2u7T6pEQoFalVuLjWIfCsWIvJV/+pjIxeqGgDsgfaWsxAZGYyLVXEkn6to
H9iY1G3e4GfGvUYgUDmSP6wTxTZ/fwMCc/MGiq7e5dIwrmd5ORq4pP5Ut8im9kUN
iW59zsfUJQU3rW86axeHR1xPNwXJOBXoh3ETKLg1tkjGw9iLwV2ZD920Pr73lMIy
KZxwOtSA2IFbTyK6reMwP6mj2k/ZQL0G7EGvlhVLSsD8GWqW1Efmvtb8IN66+yCY
JCvJPsxMJ/2bSNdrw/FGYKgezR44hiCJz3AbpT5MmjJ6BCzAGU3o5earTUGhyVAp
aDLl4YabJiBJlliPi/rOgM7JLifwHk7cx20OcvH+0PMuoTpM+n1PfEqbzy6KnMjo
7l+CEDr4dD8vKeVJNQH1KUDAqCzPMNDPdiVPL4X7vMoM5I4k4CtAwQqB2eKVGu33
wHhQ6pkwzxX5H2B9IsXg5Dyk74TJcftgX4TWNcrYvHOpB6f1ildM8x6E9j5EZezh
0LSG06nXIoinf5cn5fHl4qIVmzIH8swbVcbPy4iEcAR1vdO1ZciB4G020p6Tp8ij
/8GAhltHSYwuVy0zg7WHYd0xHg/rzluClv7Nxwnc9RuuSI4DGdKu56WBsI9CniRb
vHpRFBC9ZJtyCkQcNLSSSvJhmFKL0cWEl+p03a1hYar+42awAWQ0L1CqpogWYays
QkiZdqViHaxFykhHh4/cvNvzHbvqDNLax7m2Vf+Eq39Hnb8A3VIwUDARJMkqcRjl
O+i46ZhKsLVgXUjmdf31EFk8QDkU9RQD1mGNM2a0jaUQImDEsYQs3QxRv0CgOj86
Tjck/sYYEVpbKQzxxvewR5RKLe8GO8EEfF6OHp4L41k7rWyjjkjtnVkGSlD0gx34
VlcqkuPaNMdcgSFmfdKCbHWyGpgUwKLkLc0jrEJNadtd0UNBVP+5qaN1g175SeYh
7NOLMvg2BC6GhQcldYqefEeOtJdhwY4ZKLGBHPvOpZh0ep0qwkk45SxBWKA2VUFb
IHH/4QJbHcUQe+k2w4Zj99JGI03h0DzFoOyeuuX9gLq18zQAGliedsJ4c38HBywY
dPUyGqoc2lx6bqgRPUHPce4SN52she591UppPGb/eFMdJXW9pxNBdlOnsAuD9Ow1
CEJuxJ2afDDAeSM5URq4qmB0ZLJVT3Wm6OpEpZ9Ybm+YWSxOAuzSdGzDt3jxYChW
GxNtszeP0+eHbWUoz20UUUeBfu4xPjLf8dTu/SEQoCB3fUkPwyZWx65KWHmQMgm1
1FumAf+2F6mZwyl9Z1MraaJ0ubJsrDucAMI5OgZcsgxTarOKZptlryIc4ndxjeNo
UfnDxbrpFXzKJynMcPN9pAKmUhnyM4r6rCujJI8VhPaY+Usvm04UOzC46t7I39XY
+tyow7oIIcHd6753OfdRcnt/8cNKHgHFyjocrNVw577HThZSFazLx5pIUmof0zqT
4EkuAWTgWcw2j9ikysrR1E39SY6P5h/CTvSQV0oggcI7SQb1i2zQikf111/sIwGz
ddKMZ6mS7Klva6hpuy501Xkf1jDMDULdl+yGKNzqsJ+zpZnSx/RFjRFWk2E9iV5i
CaF3I6NjUH8Ma6GmVE6hiOP+zKusW29i4woEYmGClv1NPWQejPA3jb57V48j9Y5f
kKLOu0QBroDXRmXAZmvLjg57CEhXrI7RoK/b5cde4gHde+AO6jVpI/HQ3m50N8Ab
EUxmOAdIprnURBRZPdjucv30YIEe0OsFuKGNAU6m9Ustb9oXz4QLAivSbJtt38Jo
5y2f8c9z7r3WQ38ad70FfNiAucsCcSkZHRatAK1AQAEOIGjCLXWkgRnhZ5OUHKq1
puaJ96Lt7gogcBlKQPzEnk5RO7nqmqr+VBw0KIUI85UUeqyxnd3/10snn+fcI8qI
Hwu1HF0SFLGVJMfyseVBEJIs/nDCanGW1FZFtMsQGeVyNt8YQRZohU3eQDeMnOCM
mNnczoVEKXHOuXDZ6mKtmHVjkJlIolv8ZI55IoOKZb4kfZECMX3ZjbimaegXagpT
9uLkNEvOYgVb4wOuOMMBmljO+EUaYizjRTYYWlqCATq/NnJC5ktUoUWbnycyfnZL
8U0PyXtpRPBdrMu9r4qCsNqZD4dkD3ESYkxEsRrMdMefZSz4oqg03BCpVDq+2U3n
aShUIEpguTEdZG4cZ8fxJRWAkK2NcyUpdl+MJz/uOyl0gRCfJ80D1Vr7+8W0MWtt
UV7QGbJMtOqdkO3w/nWxPaqX8pf2sm5B/C6Gn8w4j1GoO6DHHYWJ12ul600ApNEh
/iHcUBslYb63ycu5Gp94Co3TitwOXJPx6FQAMdAZsUZzZHHLvuHWdfUOaPDGaOKj
Z17/vaGl0VBp24DxV6t/jb807BX8iASi7vLfimBmQZwcIzJMrYsJmfY1MY1G81v2
cM4NkZbwm8JTIXEoUYtGbPVxHHiSg8w50Yzv4e6O4RnbvlxbQzherm90cAbcPGPz
sS0TRlGyFrPLmOkIdoNdI+v0lu/zdRNViGLuKDQhWk7qV0Lzm1kapRKfNjLx4tYt
C2PCPgxrCCe9RfeYPusmKh5FhjAScwgfVZkV6NJv+vKDYwSR15NF5C7tYs7oKkPc
LZKxEiX4ZfiV9P/SU79xJVyf3J8XraQRujocwLm7OMIgY05IQX1IcRnKiWmKy8gy
TKDjrumUWX1GX0baYFc8B1fEe2g8FipGT01jREBwQcZHiCo63/wgrVFesEj1o+wd
DuZHe6ahGmDVGFuqo1O37T3TKZieIRZdmFGEuHFQcx/RVAYGibqeoq5C64p6d9HQ
VoS6B5Fclduv+VR8dIvx0k1/4c2faAqfu0wmuO57bblkA0yRl7snuvCGcmTlUfoG
qzQu3+37BC0/CL1xAyFaNqwnNzHjPu5ax2QXGhuUxFBkTjThCmKFUxbN2BS/IFlC
9s2D3DNKey3LVv7gB8k5bGzECgL+cxR01b/pG1zBkEgzZzcETHHOFo77ri75B1Cr
QZflMTknhLeJXiT6yhnRJP5+C0AdKC/NqPGsZI1raw3b7GnvFhzIquiyUb0BCGkk
S5lG7kI7c/C/s4FRLjuhisdr6hyWWTq8OwocWv/Z9jfxQo+U7A33PxEAhhziL3g2
3qw1CVtLNhi6CIiI1dmDN0TW3WBwQeRDdtkcel0UeOwhPnMmCjy2DpgYXTdVKUy4
42AysvjtInBbSUmsYi1Dbfu0ejMYiPob1/NQJ/+BjUzOx+KPr06aYwNHzbkuq8hF
WR8sbz6xNJDlov6ifC9g/qaA1ef6+P7eCwMru1JI4oBW9YSwSzn9HCeMWv9RdTI4
RDBuNckWlBLx49/YKZcLZ30wjkvNCo5Wd0RiU4VqmalCMSShTq1GFeHsaY7r6koV
nCG3P3xY1z91nycD7+HNGvIEc9vuiBB5IMz/J/DTa2nocTdxeVY1c7zTy2IEjT5x
d7fsgVpHjFhTD7xyhqobMLfhlPi3bNxz/M5X8cyfIOTeHXyrKjE2bre9TIzKOv3G
KUnjZ/B53Qqs0LCuASGzprqtbNEmq45mEodTi+eXAxdbJTRj0lM27NBZMN6ebeTv
0rOkNCVd3z7eMmUFGwV4kEvkrf+tUKTeaMamKz73r4dc431fOm2+AmHMak9qJh6R
1oqhFGsyjuxcueiulXLbQPd2jjMKgY+spObW5nrD68hEOA2k9ixpjXypUzqcebcN
Gn7e+bHvsHBtQbrn+95a5YlQpNlaZQtEkdVBV3gI8IpvNYKmbMQ5C971jSkRj8Ff
12QnckrTscudT2Z1Ujzf6E4wR8bqiPMlLyfcqva/loj40+vns7MvN0iM3QLlWq9y
YgukQUOkTuMHNHq+FV8l5Ss7m915l+UGxcuWyYguBeSVw82MHyGexJlrzx6I90pi
KZCFEcEVLcJ4jTUjPtc9wRvMczh1XiMwFHmaWd2jpz/nU4KmpLaiXNptHbOR8osv
53e8KdTeObTCcppIsInpdh4DSdlgEwoLpOly04zT/kfq3VZlfo8ykYqEoDIQ4CIT
09pqUEtowu58cjJ9LCpB6mp8M8Y0aaCb2JxRlvfDvviiqHoG1QDZgf5i6vBbQZsS
GtKrsqlKVGLSVQhiNxVpAArGhvPNhulNiW8yORluOHdvdgU9g4yUzIgHX4aHtGFG
sfbqzZMHpJIcSeWa+S3N0g72Ox1h4WaAU65dwswZKtv8MA+PHsTJKNL2ivcQ/LqB
N53Nwx7NVTwZorm5NHW8WzA9i9Awq7S6TESOnGOaHQ+1aqPcIT8KThNmfMMCKSVq
RDKaaCPig7kDKcnvsSf/iBwE482IZhj04y/EQQUdBkJ8tWohwp1/35f3yOeOrAoF
+ongRB5ALKI6nA8c9qP58ZbtiiBBVVsX6Ywek1zzyxvSZy3yToll6U8kXriXgE2S
alH4CYxYVsH/K32utzqERGua9BT/IiR1+pE3X3KF6m2xC3zkJz+cBKpZMBM/ZZK1
RR8v1GGk42ZwzQ4l8bhSg0zqmSTky8Yx7ih+4AEi9lWjOmk2OJf/7niPdsRWsv+1
6IpAUEY55kcBMvPCCf5UCSShx8nwjzJDSXsb8lUMeVprFfkk/ZYSvL9G6iF6G3kM
s+gNFOTQdsH5ztCTU+AuBWFwPOG8duap1QfgyDu+2GVMGQ7LwelBR/I39VSU8wIC
3paHDYnaZs+GG2i6HovGXHhm59/UdjcxbDCrVYzFPgcXeb17CD+iDm4QPKPP6jIC
81D1RQ4Q0W963AExBQF2a9C4z9H8kdY0wZSqDNN+rKGE1/62YMggEc45NyzubYo4
4MyHWHjB6a3051F02NX8W6arUFJjtGKRzklKjaouCk9id5RAg09Zc/+LkR1vWBbm
FoIhcwaSvvHxiaZdbWsohfiaRSXx+1saDD8Til+pXTlrKV6zaRBpOnSPRIxO4nq+
6ZpK0kIUPFCcTl2cyyb/Oa2kie1Fv41wj1zSW7T5SZrfq8bOFMlNXoH3hYQH4AJM
3030hcDFE1iueXH2oLUnNqLD0PnDvDXpjxosgSvaAqiamN8Omm/2idrUHwjLg9bG
lVCUKBnHrD8U2+V67m4JRcHcMRwIW7E6wnHHY2GxyIvpbdJEyWAGb8xQY3squ5Sk
3f9QH/jIY4DQCdFVRqsK9zWMMn6w9xs/o4ftf5dLBE7p1hN8X2sCVHTLMgr2q3/e
P8Zooh4JhU4XW8lBzXnZ4xsBk4RS2a9rCvJ+2o3Ic4gYmbjl5VW/3E/6WVlp2c8a
nIY214eKe2QGaM32xuZT3x3p82buEDafh0B5udu1y723j2rvpCg2hiqIiiy4q7PM
Z9VW/ER3UdRm4BJv7dznADOFtvxV3z/F7FX1G85Ti+IkMxjSMmRUPqjg6HrZswBR
Z+7I3EjZctcoBeWl1O9Lnas2UUhsnjPDXkSKpQwsftmujzu30xzCt3HZaWvkyP2J
Q5Md0BmfBH7eoz5f93yoxUrHF3HzcJA4bSI0CclzdSAGJEWgr71LqcdeXiwyCpkI
YxJ5/wU4U6FSa9mjiUtLQ//R55WlnC7IUfkOPwNLYt92iqfj/uaYxuS9qEUM0CjA
U+y+Ny+pxbrUgQ0nk6rPKYYHa8Wec4YkfOV2GY9lEZ+NAE74Zd7/fHVhkwIBb+Q3
YtKC79ffMR7JxZIQsPWl9ZRml5e3MgpznMXFpgJ1zm0QC1wX3baJ/aIWS0D6AJa/
uRbg4NDTG8SyGUEnbqzjbL5wN3UIVCyhaB3eWx1HAOq1GsURMOAuOIgqY7OXnrZy
4ryD6NSl2idpBpXzytFIWFwf8OKw3onKKKpla1A/7t44lGdQkIgqREnRRYY/A6b3
HnmC3Fxr7Emg4bHTC3Okx5ogZeM4FpjWuFr29KA3DmTXl7wbFMbyrwkJf99vQ7My
a7bSbl0FwkZ3hKkPJwEgg601sVGN28PNKn+TYSGKXq44nh4+zLEJg+4IOjDHrzfc
LPT/g/yoC/pway3oQLSWy2m6IvbJQdc3zwP72q/0l6ld20F+nHyXVZSK6dT9vbzi
TB/0l0kFdTsM7p7y8frmR1vHNkUKT4yMAXk75dGI1vCnyvQyBHNaquUlJmB/OPI6
5vhfkj7GQguHVpPewM5OTNT5uHPpiYWodSNkdrnG0ZMAyA8vxN6mKw2NghUV981s
qWEXZ64rxHjiKgEKkHlr4mEGeGrvnFGd6SRK5B7LQtfXmwDGGu6lISgTjyhxYYio
lms8U0CLhD75o9KR4Gca96nbJ9Vju+Qm99pWexS7yv8Nqm6LS1PlhEyLtEH0di/F
zo2P9Oj+NAzZVGDNx8Fm5537xBeCz3LgcFCNiyl1maoWkOWFsLSbAKu/pe9G/Sge
Wfu7OHANpJaV0f0JoMhIeag+ogvCijlMcwqLzcJc9GiO52DAlAWAfYS8SHkD/eIs
msJT5TsrWcrHf/xdJ6CPgFXHgq7V92CVvIP2a70T8pssijSxJGjXris6k4F9rqrK
KDYhAoYYToLjipD8EJ+k5rSxXLt+aeQxmRszHIiuDLzC9l8t+VKn5xfObC/DNfoI
VV0zMyCTwRgnqNnh3bPC0NyxazQzlnh1bnip+8bOBms7UA9FwYUxWYXW0vswQTi2
PkYpnNaLET/sRJdDSr0j2GeD+g/RDZhiuAe/jD/6v7h69ImbW+BfP2ABjj3tHRHp
QOA5bmkr5j7x/G0M6mJOHAgMQEoM84IYjfxgTIaeT3cQAcgn+ABl4s5FdgONgKad
KtPQ8QM0BIjivFiPJPazwnC0wbP0o+7zqHrZqHC12HqoPaUWU90l3nXyaEaxpMZL
Y5dQ9H7yCgcwioBrbZ7DaEXva2cuFhvoAubZTSomt8LgeF6ybvXGiYUPK51/kBo6
sapVsRMNUfzSYW3q5g2K5l78I0hM/kXD9vweZHIYepDBB2McmKeiYW5qC1H4Ge/7
IOUyfu7+LAy+hfiriLJQQVAOWKygF/LAddo/cM85HObgnms86rjc78hUIuRVekbI
JuVuU7anqsHgtCyiWDGCMp13FP2jkUZj0jurx1s6jlmhRXo60EEjQpV3FCXTJCt2
EVXQhhyl53tO5ij24Q/tCpZsgoVlDtRqLEOpYoK4bLIcFwbWFW9X+XOhn9k44BY+
LH4KGYDA1LnR9A7v6uP6oCTHIzDloj3a4q5HEw+XIlkdpy7REHcuI+3JWnTA0xzS
Qc//qMjh/YReW1d65BUbvLuPXyCTafACjsbKU/TJaFTIUK6LXTbuFV73bjgCrjCa
x9b2hm8e7tzgzRlZuWMJkHoDpTkEQTUDLgFhxRYOl+4cbBSfaxujOUBzm83odMRM
WFiJL9Pn7JQv7uRbftYgM1VU1VbDWu6z5xQKHmep1+kwPi7TNu0kS5LcKYQLf9VC
Ol8876TKdaL2IJYscU2d8IpGAN5fsjE1nqhiUCfv5OfXKs74Vm4HN7o0Katterna
Q9Ws3VPosKSyADOrPSIIk69D3Vmlaub20is1O8IEmWB0g4WrL5mZ54tiVnDKuqEC
C00UTTT+RAQ4nHLjJ8U+tTfDGdlCIp9ZEWj2t5Ws9kJX9sMtIMevEA3CHUKSONcY
Xw1NrnSzSjtW1HJAWB2qvgD+Kw/2OiKQQuFZP8iS0Ez2SLYz5vKGe53RWCLjFfHL
FOqwPwctJVDBVtG5S55bONvsvRQHzOLoogmppfnM7cSM5e4YeiivY2x3Ma/6jHlw
2r2zWLoxPku+cY1RkS1CKMZOlAtj2LQPbzO1t+VQKWDN1zqwn2+z+A8t0ERyT0rJ
7QD2JVE1HbxI1+oEGBI+essZ6BoAikzn4iEJtXNazvut4mBLrdRPthP62KDrcIYH
PARgJSWg1Zv5jgLth+p/onl4u3z7/U2cBg3R0GwaNYr7G38khJKa1ixx92yKsdw0
Yt0ZQElUNRlyqD0QU6dRtZ7cxCM1KZPvUv8NYwzB2h9c2tyRs6HpUbqTk+8xFGd6
wC4VdwpaZb6pM90IoztGZ7cAlOavaOs0jtCtlDasfk1ZBvawbluGTs9Wk7+NvoKV
ZGfAfcPpZ/vqYAi8ws2XSODL5N6hyife96QIZ3FDsiqMg5CBOsiU41qjdKmuVM+/
+OcN4yvLRja5JwRGCbh3UY7DxizukmGsW8R04TzX3p93SNRJSC0nqO9Iu4w4HUXI
5ubuvtJKre/Zon5k88Dq+vORB+Sv0/Dh/UCcR6BjimP8UrV1IVogT+8D8o/R1Hjo
FXdb77uIW4qI44zaV4LYcsHDEzCa8yldXZ6xtHnKkopnm078wordAGASYazV3AuS
D51qJsWm0DdX6gqYm37AT3UdufQ9KENrDMiZUZVbjmn05VydNpwFRNl8yGShKU1a
2RrLLEHgj3e9WMvm8ECAjxQREFhNBf5v5qDpykqTjPb3c0Wbfd12rPkjAaJ5f2Qb
73thZbBeBYRIOHRa8r5k6PjL7eRoaCEC4Tzt7F1erGR14m+mvkkzFOhxbGK30tRl
FYys8LpUaAciY4/w5eP2xYy3n0rACtVFali/teqqp8xZmktnDpwVXIBEvSKzP0AE
8sj1TLelbXyWsGwA74fg+VYeV+w5ATtQDUsvaAZ/T0l2DRcAhwkj7mD42VlQZVN5
sGCJGEpF6pI8s7kKiaaIODSmqin0lNnvAihTCUHioEpHLcYUEUJSkaVvJzxRchVX
VBtUD0a/I5YeqDGj6Q1lJArxgUJmfabhPEsDVaq3lMUVZeLQZW3WUbRI1b3QHlRR
tGxfSYeIkVzGmBGsYvNNJfMxGeQ5BAXtxj82XHM602c09m9IiXYGojxGI6W3OnCE
JstBEUQ+nZ+uo6ZKRA147gdxMB7wU2J56BgHHhClpe2pckNFw7fSuJ00uua64AFs
Rvi4kjB/qXffR2RKWNpeDaV5uU86BO7QFvX1HaBaZJCBw3z/5Vds8PV42Y8Sqvmq
/pfwosf4t5KPQcQjuhLmpUa8/1VygNmYViKWt8/aNhJeo5W+xO17B7Nc07HHHOYY
jRtN90nHfsBVxFL8cHDsoW+QLgi70dEe8kFEbva6iuXi8zfsauoW9sG/Ub6MMoaQ
usL4JONAo09aG22pdsNTCQWb/YrG5+c1tzntGHz+Yi34uByzEMkXdDREDI6TIfeB
QA7re1/7DzTs01DZd4yUSeBTLiB2WBm29sfNCjxnp6MGhbuwgoltrvZ5U6C+XbEf
jCmG8xA8PzmLGoQ/b6j7NRBvA06lqm1PFyYrr8rAmcfePRx7wf3UDB5JGty0hlKn
aFIdIpdA3I9H7fT11GyO/F+0Ma9J4pqaFUFz68DA2QaJ3BW/Flt/oqf+/nPGYDxH
n5NzPU1/NqTDQr7iuLLDbm1c2Uo8QJAzpdUbpTRm1+Gk3SF8lYF7VgBfgVJePRmN
7Ofi6IiijoWWWS28yMiB3m/8YlZEGyHEDgVdVpB4Fv63D/nH/3O6AMJnwICr7/TR
EaqPLS/Ra6aA8IRrBP2aH/4yEdgb6C1hhJJTCS0/Bwdk0ChP2WZSNqqn8hGyJD5b
/D2Vr27btqrvguNsI0ueGPzqbLWTQaun5apSToEw8DiDDDxJqh0C9XiSFnz19v12
yuFgRYc5sCK6r8UYX6nxjFY3uzhYBSAbh3dIrvOKHxS1fAeRH6C06COolYdbUc3P
z0LgjOxsTEJtrgHhS5YThnVociN29UYczJNFOvtflWSRZ420BEi4b7V+NGWF4ZyI
ZQO1SmLjykFHe5PHKHM5NRpJQcdOEMpvH4aAsTcOeOkbfjEjNeZQS9ZKR+RwYlpH
xFZl5x8Mnbr+6wU6AohIw2r4uhTV2pFv8+7mEb6PC5BCSmqu5Q3tjNLu4uZsQull
JFZx7iGx9DRF8XC6Buelw3CbttdG0OnHC7wxECHvV4wQ+YNmqEdxRsAE+TT6Geix
G1r5Ahxu4QEvkZoHS8PyxK35/gvmWEs7k3VdzBFLccVVsMvR2am6h7CJwFHvctuG
wPBpbaEPYUl+jiXN8mjfQYC70mXo2Fih54bX2Pwt5K99uimaYgj9Wr+D/iHLDMCb
SP2hAgEP6HjVNXF8wVB+Gzah5mPGnA+lBPkgUidyhe4uKWBTWVoOf/KoUX30a06T
LG+hACNsUZqb9eNwQKX07K7M18Py2GwqVFX7TPZAXU0sj/52I6dhNodwuFYmefyg
7IYExPLb13YdAmhdOHg9/ADQ42oJ4cZq4rYCHc/dbThVPGYHLeyFEz54dACwQeRL
LVrwJM8ZEjVeFeLGZr8myjeFFOWi+VTEs7AdwJxbohc2k9jXZUZ/9ke0TFd766sM
4u1EgvQS/xf3NAwc889O/3/HotlyGbseibaoYlsfKAeLupgjGOfBIzwJ+v7rK2pV
3L0A8x/NLd738ca5oZtOJiD2Bvp23MvAjk7+zgIF+xBIMvF++a9amFpM/jO09qb1
x7VyKPbucQOairyjbBPd+L8zUqoMrJfn+ULEDlMhMz4LpiNC4krwgrCORn6eKXPg
eb+1DbI7A+omB0VVIQpRSaVz6EltxWmpzCkOPkwYJSZEBEBCgbCTvFTf7gCxgTwc
kyMR8Cp8Od5dJJOk1s6iT6/OLBwouaX6nGGGhvt4dNTLDX8c+O7qT3/8iTvTD2/F
DORFCLOlHclFtNbR7DILSOxWNKaXMdklE8XZu4TeRSVOoXWS50hXl05JeXyNxLS6
kgUuvS9RnHjKTjlHFZyp6Dt6FoPwqAvZG5Q9l8Kj/ZD8zcwZInuBZOwtGC13Fm8i
Fpgm7FhfpMpzW8+5pCeKTF5mQtygqdHbPaR3G6V9F/tKpD0b5I8VAEP5T9Gz7k7n
AFoTLIX3Up8M5oTahOYLCsd6aeisgRGgF+dHKOZEVTqVSHMY13bt0BW4uB2UOW3q
m5jmD9tlA51b+fcUJEY1zH0hUt7SDLLCGZcrHcaC6X7MvZBwyuuSN+hr0C4Jx6kJ
oROlfDtJV7DK0xDXqkvzQSm50gjYAdDgX7QpcYmvl9ZLEoInCB4f0gWx2UmjP3wN
eiz4nW/MJL34KOl6lBcrkQUlfXeyOTsz7THHQFZYLNH1tjwg43v2K7Ua4ZmaKsN3
JrhsJeEanJhE2mRaCSYxAYHWvjEggO8NTLWXMFK5JAMXwWeLmptdFdL+Ae+/vEnZ
dadFdCXDmFEMgEnxQLCh9iyWUFxA3vD1V3sMqyAiEX3uzIxFOg47I/bnHapauGwC
7R+otURsgxTi9ufhWr8eeiBJUJVU2kkXXW/RhbOufl8+KDPXZSBFUB5EWoKmJCc/
fhATqUtbOl2uAKcnxMhK1rzUV/Dcf/B2LeMHhSm0IKwH6HkHNLUo5SOqtma4MAMd
B2NHzo2UFZUzW+QWDs4aVCIenBLdfRiOdNaVwj5qAqx6TBFVBQvGM1CGvUcLS6/U
CVLqkhAnX5mPoEi5p0yhDO5xYfSGcVU6rp1OiiUpKIIXZsbXq47IZqOLyevQqaov
D9nTMLgvf6Q95SkJWALrwFRm03/Qtl9FoCipVs88Rlle1GSan54IDxki9xTSo+cI
NmjzMeFHL92KjRk/nV+NHPwA7m5IyKENAYo/u97G36GpEX/XJPhqZCTSst8dyWWW
UFuKk9MXgVq/ar5BlA8B/UnFcpdxZdhP/SfwB1tmaZyDhUrGNX/Hs1sIwMgyUG9H
DihfZ/GcslVJlciLSdn3+CuvG4qQxBEqEKa2EcgdlefHBHM11UhjcGiUJuhtTn2q
evg2H2jF3gBPMwzNDQwHoElSFSaX0+FSE2ySmeNi/IKPsAxVNX9xC6MqLf8H9Nu0
+eCuxXwpxZXMA3k3OaVzbrgxKHwB+eG/Peau+ME0Z9CPGHSv8Hev/o52YgErl6AE
JbOcZnoIn4AV1b2KhZhKjlix9BFq1MSmkKGTjUIQcJriw43gmQf9cHZvgNXux+R0
TV07FmCyeVeRAWP845vlObuQnOn7FykQjuxIFQBDKJyFscogLxG5NnmgzhyiOI8X
JHgEH1QZJSHsQjx3xcuN3FT7EGBi53AcJGOTyjjwwpdahF70mtvvpn3T4FD418YZ
SKlsoJZZjoE0RnkohDL0xDTlxpnxoEc7QXsJPVX5lse2Sj4Bp+ky3c4uXYkzKL9g
txY/4FkFu7v6L10s/p5tk+gyiz9XmN+q3NLU3A4EmmxKkgUtVvy8SHhYy44wpDjL
w98GQyHNCRuCJaD7HmujPZDMYO6qBbaXYWyQPsWJhfWDAySKMI0z6JQa61NmM4Xy
Z8roTPizqubL8qxWFrq7UO9k2XdkZUXB5F3wDYLzpLrUyitEn7Hz/cZdTja8Rqau
T5X5mKzzjCbUmL+5ww+/mpKg+0qgOiq7wjfvWAgsb+TkANMJArcBw/k7Uzz0TWd0
6iQPXsu/2apNLzcVKdsvmn7dbSrJDz1lDuronZN4uEOOFwwlNzzgXGkw+epXDOPi
hmb+5fIHIGjvTqc5h52PSQ4DGPoM0HP7SWIbyFHMf82l/CGsw2xaVydmVaHEExxf
ItmEV9uBQMAVHzYXYfhr/8eRiSsSFk7hg2IelGYfeNtyTdkbQimqu90hp8gGalVa
2Z0TgW31+mN0i1J9aCLKBdEeBvr7pvnpJoUkN4LJmgUSxromaUIktHGTgsx17oq3
v1euaK014AFXYKdjjV30cCK1fntBFjzaotEEQNtnvdozRweF2j43wwOGjdWCjdwJ
QKS9CBsMe3TskuhZaOEzmfwzBndpSK4Mqjh2k0HrKu2d/6KI7LV+AOA3t6cMazTa
HAnLY+jEqGwIeLFVBkOdccUMSV623lqMuyl1Udy/Lol0IRUvm1JkVEb6YPv8LKgQ
8wLW02+dkJ2Ugddbtc0XnH5zuhgpnHcxxfugg8OtCK3cWwLc2o2jhKiNFychyOai
XDefMtyqTtXNXsURHdeIWly0UmmsuvuuANLVJjqn/dc1ktR+i12uQ5Kc5FSY7Djh
yLnVgzPfP0bQ8Jl1bAy5rcPMI1T5OIUhdbfR6DMa3gZgPsCwYT/G2JTsTuQqI+cm
JqqDqs/c0phuK4e78ElYiYoY1xKDaOw3CK6drnLm/DigerRPEp+dgP1dBkqZsHoc
u4eVF4p9DyrGBAsJIF0zte7TFmLbpTwpWRpqJdoalY2u3Yq4ZLCdzR66awHZqO7p
+0rH9f3G9MF3WqGFOXLLsZmnGqMowe8YnT/Xb8TTLRYk3BbLTi1eUKveeij91K6a
ouNcLmXEV83MEG9PEvQB6SlU6RSWHirwSyFOV22oBafEOdGw+XVD2yOX7tfMksgk
u5E02uhFzrsAIibdzhaWl9By+kVqVpXhGb4BabFchpABRpVIYyl31zLIDaYxj27H
/9KXEbODm48JxSoyx5Uw+VGGoRLU/eIJjwOp1PMwK9DqKMUoqeV4I6M4Jovuoshq
0nlbxeix9uY7mwWic768aqiDJ3KumQNwUNsBv3t5thuxiMFzFA4mVEn+q8Vh9rKQ
QsvX3u/qq3CY4k9ibBxxkhhpEK6CGjMnROnI0SMVJ3AIZXmX9+lS9Umf3P23DpuS
Q3HcpIu6IvDbPeftfOCw08XJE2NXW7RWav8cqRkPFzB+aYkhN9RG672ik4xOjU0v
LiSMU9u/60tEVeFZ4YPhD6nedVokaAX3moaqxwFct2ymoYVebtR/259mSLF6Gdd0
UKBOPvGUT86/pMsQzjmFlufr+6tNcsbUnZzV8eeRPV6mS7tG5msmtKYSO8OdBHWr
wNNenI2A1fg+9gU62w4QybFDzNbFjP2goAJseq0Geq8Pf3UAc0yDaGgE/P9GGjxL
b8bB/JJn0CE6mfMT7BJGqIfWE8ANjmVLdm9PbROgJ9UjS0HhiriKkgcKMX4xd45V
QH6fVOpXLAAu/gMtMQlQcciCYd5a77dZyBJpoUo9q+QXKBSPikwFzXQDoSvBOE+3
rgeVKVevl33+caXoJvQO08wSYcum1AKi+YSbr9cVYmVXT196nYKatur2yk0fZPpR
tBi/d9jj99hsgKTUc2qkYWIstbBJDh9ZvZjBX5Mra0vVwdxY1PqdghfI7+OK1xX4
Wmfe92Cj4ba3DudcbOztw/VGD2pfYTNpMsyDMF35lj/7L1ksw0Q0ZEkMblnx8oiR
FzWSzSuQMwG5DbQEpJTnhF1yASf/SgZmGA+s6RBZQQqA72hxddFJR6x1tiEr8FKa
GuxE2q7orlD0l6tXHsPwJpktnAwnijnzqezVYasPPnSaeIeI9EZJN/yL8L4/79Ul
hLK19AmhA7VSYqiWEVEKB0mFJVo+FY9z5FlSGmNAGApGoUPEx/vmUwSFTSjU9U+b
93/72ZYcOmIBnVv23Bx2pnjR3BQMQJ8Blp2XItusKig4kWicwZbi7DGi9BJEyz8q
L1V2NGGDs6WvqHn9smeGnsozGr+v4yuBgPGEtMZgb+BXXN6hZrD8KinCP5o4ANE/
rGZIlj4+KP6WdIbllVhA3NPOp9mbaDRMXyakd70JVSJVLGvQ+yplQVUJhMo5E3rs
FwN1pjy4C48hv1pP5O8Po8HcUvoZt9lCuBX0CJTe9SzFMIwrdBcS/1ftLU/gbHrA
tCyyl9dUcjjAufLVDEthTI5dHHnHrIPkO5GGI4XlraE1St8vL+V2vCzSqCW1kYo9
QgeMUrqacfSb6bWZjSq5V/1Gh8fQiU5xYuQN/3T1FP8CKc1488KiuE8rZSX4pdzC
7WYoknACCu1qRa3tqnx92T9Blr1JKj/m4AXjVFKdxcBUdJWSjB5bURSLmWgICYSY
+PpJ+84jlJYsLBlly44qKt4M1JR5jxJ6mcK+67UZFc22Xw1V7Vuue4UzxNQx+n2i
MOT2Yu3w/UM5DBiqo6oBbXf3EBStMJP68Yg37imNVDkgSjVt3x3kktqKXEJSCJiA
PO3Q7tU7/Q/Y/apL5CLM8USlleON79OpTGoa3QQv9yhEpWpccnyG84r6Hrqssl6F
8HotDMDUDKIdiORaslbE0CRghJ4zR888SGwCcIgTXM2h7EhZ8Ndn9DFimPMRAEpr
GNYDAXPsa4a6okE1uAPYyYazgYBNDlQH4mHYHzjYvM1ZCZm/nEb2ozKZ6nFBqxbD
mGZ22bSsP7rTrgSH6YqLFu5D0Bwzkv5jZypQOPQlcXN0CqNkyt6GxKx0bVW8wxGJ
I6aKJrkv3GHFNWrfhaVTaOBg0rNOg+iLQrwMbhnQT/3r9u0tziFgFCDCwZSKq2E0
nuvXg2GHzOsEUssBOwHjhZhbq0bdCUN3gVR4Db5/H0EqMusAiy7KUx3jXAwonBKh
N0hO77kIh+kINMFiZIcD6EBXadpU49cs/rUf2HDuJfEnFTWBDyY4aEQjyaRQoWVR
MatMIxTAhb7qNeiIZHIJ20qtgQmTFt4kj0EDEm3mwYSnb5EI67HHeufL0eP8TF1S
5T0TK8HIVe5tWfSdV9RgfvYIND2RW9YZt6UxVhf/ADXUrTWVpOHsa+MQ1BuxdpqY
LZikQCt4O1fgzNfcC1doKkkgmaljO4iHf1/OhJPmbgY1yxy/3khImkqhepdTZ0rO
iSKRi+DI/1/UrxE5vp3sjppGNYE75KxuG2D9jAusQFDiTxhQHNcbUM2se9j2EeET
4NHxt5QkuAPtKTNJJIgFf8mI4FgIGuA0xci4tamfawfwcDuMxwBUrLob9nKHnxqA
BkYilNuwXubcCNCEiUOkGDvqAvaYOh+XCdgMyYt35jbZiJNzrCZGEPZyNV5MX7Fw
OFDaS3fD0JR8iUIXj2tICLW2vQKnz0ZNOBOMRJtNKjnq9AfYNCuqJNq6KecvkX4O
rxlTri7RW/+2n4AYetrRsugDPr8HcEXN8+s2iQ8fplBTDM4B5B/c8XFbk6hJ1exR
6+JA5fUt4+fOrV2R6W/wGFGgMk26/L/reCFmDdvhZt0/d6Ptu+4XdhVOMd1GoEuo
NSoPQbLXKBW6Wzer3y9QwATRXyT5nxL0X8tFrYvw+z8JCrPAAsIMSTHl1p/lE/l9
P9pLQVExTIq/0BaKSzvkMq36ePweEQUD6BO9OU1J4q0dX2hylAB0RdGRFL5aDcsK
7MM109RcpFZa8bGvhhOBv+XCE8ffaLHbE2TURAVUTjJdlQaKDYLtJnFH3ti0o2Gj
jKyz3AIGsxiY86okqCYu4zD1YPji8KPGwFCI209xCaFu3DRtgoqDBrwH+DGVXlDV
oeBylF1+YS1REnxQ9T5+fxfINZ2RA82FKk6LafYvWVjHA4wMls/UtkcDehqvWp2/
/hJ6PbxkS0DSDYokfRYsf99N85xqghRDVU99/DnMyHpePy40UkwqbnIxEHWd67yM
+j4JjGtyBI/mS8C2yqDFYwL6oZ4OTZl4ZbMYplboik15W1QREt9cY0ptcScvTSvW
BTei3lrCrEZ6G7NAm28IqP2O/7SvfzpsBQbVESvA0WYSGgPnGGyrwSNoF8ZJ0pL9
1E0vaNjTV9Oe6h4wuSLZNwi9D0uqCVmxi7TYZm6YNa3zmhlgi5xY/J86jSD7+7mE
eQCI8wI3mAltY7bBs3r1HGmOaSbJ21HLUzUl14pYW56u575OT09wvh1CSjtucMiE
MjMfOIM7V3XCbDg6Ue1AA1gmd28RCa90NEmkSZXg8LK/FAsYS4N8TVJweFyXQqyC
YMFAgeZ6VrLsyLoeH8rYmzyKgXm8inMHjlWDYPnvECw3sD2OGH2BxzZpbTGkDpb9
SdN+OuKZ2WG4xMqq3nz8LAUCW3096ByBawiTqTyw/eWD0FXIBSTf6uLW0HhmPdXJ
UgJ4JkwGIQJ3AGGZUnE2HpMW6+n5UGxGL1IM6f8IbSDpb7F8zCiDTOaer+V0cvyP
cFl7YLwmZJwYHI5FdGlDQgQyG4JIb+DK1BTSR17ZLmnkqsrj7XYWurz1RahlRmxV
c3oEItRPtcorgoKFkB7DnwUxDqf9LLDQXArvahYjJU9GGwd44Q+ChFgy9CS73WVk
4piCj3UfYPLEBYXfIFAJxeLe7JGt6mo0hU9SzWAhQFv8S5Ig2FYIi7FbfcxzNXR4
MFNIDFjG6/HMEP1ShNF1bKzqJp+qwN1arbSuDoXco/dORApiQi6lFb0Q+QFoU5jZ
Nl0hJCRinGiajYGfvZ84l5CX/nIYdpj7S8cEIvUyJD1wSxEkF8vvMJsnjv2f5rk4
ggodgEqX0db7jTGICZlCm45GGeXa2IcQllYp8XNA9s7ABQBaH09fEF7GOFtqVTPb
m+lUo3rBdhV8sI+grqRMhZAAkmR8+QEBlHToxvwiNzp4mdZA8ONjMBt9+VH9f8aD
BnnfcAjvFEmVJzU5yMU5OvqMbxsTENZQOI1zbupsS+XThmZzzSRJZIirlyref91E
FT403LDHJEr/FKx8wcZwPXuct25hiW8IcWmHnjhRoR0a4RHEiZqubPzKfcag5b6Q
AxFP5JkSp8nGOX7L0zzGhHlBc8FEe/FVMGaM6dLchxP89BnldL9jbl9nfoAtP9Gl
OqtpApWJ1UwtOiQ43Qe4F4VV8OBLlVHPeQqvTooIc7B2wRC8nG5RLBPCBofiFjzE
p/FM9aKt5ZBep9Y47C22y239BPgAkroy/Os2idEX0NMgWqhI+OOHUetGIIryK8v3
2iAogEB1JO8IFtaJ47oNZqh3nJcIxci69ifUM5Zdaw9uY14ePxNqoPblSwnzlxA7
1BpTJk06qtBuxKcKW+6IF0Xe8nTJWQwTSh81WK1MIT3oBipl7C64A1QAJ5QKcexR
2Hg7eNmeFdx3uRhen7Z+deDxtok1Sm8sObMuG8UBHoU3kCq+Ssm1BryIBV+M/LYB
cAXB9TiGOO2LFT+qLhifQqiKxXDEbwh0kzryj05AP/+K0eaQddqqJrw0pjMtOio6
WBB7wxAj9LYWG97Nlv/Cq73nDyRaxqT5hpZFyzRnNms51VznIKG1fShQ/vfVt5lV
UCU1tNOuu2LeU4y4SZgrZCgOn3iU6bEokKFhaTYdcbK8efWqn5s/cctLDGmO1aOm
l1biGoh+WPxRQ3Mgz2bTQugd9CS+evpkMGaBSTty2IO4RgB3OWub8hs7VPMiFuFG
K3yCuEG1iVrjs6K9M47t+81QYg0ftt7PYIqGmyx0ktFJX9rIyogdLEmI5P/kYpKc
lILmTTml4eUrOmdHxr3s0bRPqHm6JIfrATK75n13Lm/zawuZb+85FLRRMjnYiGVy
uPofwZqWcEstlDKZdr2E1L6sQ4ZyPkvmVMnRdjjSsXm4x4ZaRENX7KKFZLiCr8uo
UFJN/k775ax9f1X/NxItlrVeWonyNoXJvOAsDpVHGv84L0Z5PcNkrfhfhRnCCf4+
qhO9c6USuSJvnmt9shIzSsj+CUfASc+RmXkTjpAAgEjzqr3VuYDE8Nypbs2Vf4sf
Guy4a6ojIrL3l3EyTMXWgZOTrUe7mOnN3dQmVuLZQWCteq8QTAzd1ZKbEPnxEbHn
70f0LGne0JSs6496QeYrqcBMrSre0kf1WL6LTv9XsCjJaf9dX/FUsP9fH7A7nAQ5
lKTu8AmtfSOEyHXJheTG3Rr6WozSd+wWpBVvzN3MDkrD/QdkGlUQ7t7nqcRK8uWr
+jAKIuwOMvSuIJn6osRT4phfe/Padx1eZOgsxCfuSt3VaIDEEGwgIqJxYo9GM9G2
+4SGEqzHCedlhCSKQrFW/17gCYL3Y/KcYDfBKi1NaFkC62KQ+JmI/o0yosec85Mh
lWC8Z0Ji9GIamtw4own6MPZ7qukdEMBMijtvfsyw6Q/puG9rW+7YzoKqT3Qj7Vd0
iXhYGjwVV+ho4XVcVkdPki2mEcwGhhUjpparOUEN8uB1KmJr3flPp3CAnx7sc2Dg
WhUpnn/uLym6WUaaSDkybIzywDdHtjKyMOHOrdmpFYxtDnF90v7k+8by+lCYqQ1V
7GeT7RNO9VOQe3GRF7Pe9/Ujid/PEykVBh7frxr00N3rH4e/sRLYBcKj6B31aQpl
a7Zxpaw2FvuLqbIRC/+9p76O9OtIFyaOL6MrsSrFDdjSwdt8RnpSZ9zHs3OYHzry
khKyMIa5CaM943MTH+XzVkxG6cRE3V0AqPruPt53/y4aSOXHYtRlBpcAqF6mR8h5
P7ZblDRJBS5Qz3jgHEURXMixKb6YehC6m4LEfO4910I5uK+62LbCT5+MHzyeP17r
CSda6mz0rzNRbYloWZ7SNuvcSq51MUC9+Fjuf+TTvymVyoH6nltAB1xW870uD7mi
vqmGNAq2Pg/P8bCY77wWnVW3QetVZOwLWVs2xW2nyF43b/p3XHVauiIn4ifG8U1J
1zwa8ic92ITlvcf8vsClyjGYHcLjT3YjNvyypI0JRfuUSoJ+1dAROA67u7kKS47p
NRGGhpJHhxu424QhC3BQIuefkMZ4LQlb6pKsdL+UaPfGKN8aQp/RGpVb6oUoAzEo
iqNddoVJhy78oxSYnEBZJMGiV/KXXl0Dj5oidt89zsg4uiO7LhOBvGAEe0VRDDt8
W6e1pZHgPL3UemxOopUbFiAvyacYRTVnh7hCd5ho44yPTI03j8J+sFvc7fNVgIsT
3F4m/rgzCaDtkA+8vaqSTEyxuYSTiuLvLrze5HTTP4r607tTj9NFoXTLbIXQCuFE
tNOzRSL9AQV8L7l9R8dV5E4nZPxDPYwtFTkMr9Fkw2dRrT8iuwU4OfPB3M3//kLa
9c0YTZ5XcVmKXtvDsCgg36ufvQ2MxJcamRJ8zCNBRIcYouvQU7bstjjnsMesgLXA
IAuAtB98GHejkvCuREceVzgrxywkqz1tnM0RbxChjr/puxYQGyha5q4AboEN60d0
DJdv4+oVLFjAC6rdJ/DKF8tATeFvGCyLQwCwO5tqvZfop+qxN38xYFlAJdaA/R8x
QJZAhzLo2x76uWLyz+acXJs/O9kLQv8WKy5YHd1ie6uHsNjakIHcZ4oLzfGfIt/4
O2DhFimFBIgw58b23sTrWHL8+EEg+CB9IO+i5DGAlsbTUU369FUpxeeGdUMlUrYh
3fCN+l7pQ9vcD7LNj+BLRUko5IAVEcr4p70GCSIP8WRptSRII3mC/mbNV6u/IWE8
qtAam6NuKU87E9luC1V/AKTFWtriEA9Tc02utYnqDDHrZ6iaQyTHB3ePKmIKiFnQ
izPFwPzIoQr4cxDZraQT/UTXXc0OemCpaCsfDBkiIRqxHTE1OKR+gTX4tKNl5gWB
rzKnTBNr+pBbo9xvq/l+ZWSGS1vVlmq5vO6v4fZK7ncjNZ2gsZjK+qVQVm7OCC6z
d0/QZrCG50u+gZLkIJ49FxMczCqmCN8Ah5ZG0Sjg1jxge3gSG1s11ANvBorEH8JD
VldOuqmnPp+FI6YQIFPSD+yPKDn7UtD/8MbHCCrCz2RErC39OPChyyF7VjBAJAJ4
z/nBz7fUT2FRuFoZ2LRtE9ha2Kl6VuU36WRyNwbUw2YaGSIznmyhlk1RUWAanBE+
yokN2VY1qsg/AGbaUCM+dkYolO5c5hUmzSOdPuqU/QQ4AYUW1F70UgZ35uYYjcxd
nQ/G0zW/WwdY70dueDMvcQoIuS9cr2HIIebjTUFF849ZMs/zgioCJGDg0/94knoD
Tz83WemjjyvL8HQlE73Ta9NVOfepS7p6Doh8weVku/K9GxbIwM4Nptq6kU6pSqgr
YWd333q78uIn8Zv4z0sYKYhtRL0cq/HowT71nYO1v7CUmf767sApHe4IcAVSmj02
VLpdwgNDICvS9XrmI6X8uMbK68BLvjzlocA5vX19a4fNL9Br67TtRfoKH06jBN3u
cNf1svz8r8rEbhwRfI61TkibihFog1P0U5iWwv+7sojX0iQ1IhLgJCSXtP3OuGrv
GslrSz7+OepKRDgVCCBSsZjtUkEefd2fUsLn2E0nNA9FwlePIP+GvjKdAhbunHBB
70GlL3E14p1KKxaCsU7F6c9Qoj41Udv7Nq9ApzCF4A3KyARQwrFpIbiThOaF7Fa0
2J+QDlwlEPxXO/VY0pIFhUyvQ0FLNHAQ2nn3I14/zEiECgvQptLEGcMrnxfgf3Ir
MbLIrm1GS3dm9P99G6VbpEVGtVhSsjQf0RmXKuHhIBJRJzZuK+afUGGt1WRFzKC7
Nolrfi1rudk7K15VfX+6u1/OjXR2QlfFIu23AADhiwl10BVOEK5kmRU3H5wNO7Qq
O7ssTAPDmndJsGi7ptbKt93qhHqDjU7b78cUzH1jFUYDJL5qr4uxnKi0xx6xdppg
CZqCuoxHL8UJ6s5ExvS71plHC1M+OvQ5SiiqBMbTNRWkI/34DfLvTdXjXSICdQ5h
5EzieSFt8B1vH6FW40o9mrY5iUE7gTzXllAy3+v+ZjFlfGAky/Y+9MODimdFOYpg
jRpBjOVXQwc8PMS1eMjN5PizUU418raZWB67afxgiQ05n5hoWmV9V5mc/1+yIZon
qhhb4QxvQAKmArfm3jEXNQNzlrN3iu7qpMgJZGbuAiz8UR9laOiwOHaef9cAbKa2
m4lrseUNa+6jrdjAfJ7eogIdIgjsTr1jRqjK5iBGWogBCaYpPaOeQd45nyTeaEKV
gKWZ1twu2IBqiGDyNgk+lK7savOXJNYwuLkQShX63rMZh4Gi7y1Oycyk+G4RhH6S
8JyImqTTlZA5kmomLefizlBECdFLowoA3PGQOrmoik5tz+IQu4fJer9uymLZUNaL
szTNjExSR6+XrgvXmqBJIn+jv8r6qCSx063vLyqW6gXtvoYBvyrsQaVjDem6mtpL
L6htXhk9BTkdLP47z+YEQwWkHeFweBOHnAuMwAfjrzq4qJ9hnczZf5pz8lkyLhOW
xpZT2SgSqaOkY/J2j9E5f79a9ryjMGg5B3SntM+e6TvxOyWs1uyBY7Vy+bsYnlUj
PeVqDmfTLUmjrsbkXQQjl/DUGyB8FiuKUEqPCG8wrbB2bjWifori3rxRmv8XWeF8
/pHsXdTMCXU1fhK6dQwTWybqf7VtWoYJXgp5J+VFHW2ZYoEj119VmA8NNz6bEG7H
ogspacXGdKRrC2NkuC1I2v9r0cReGw27odYsZNxFHd8LgJUYri2212KzUqy4nG6n
TeCoY2h5r0RPR1HapcyG01/HcAin9aqin51x7rRv+/JplhXRKh2wYXQJ8HmYlrDg
hS4ge9eSVoMQHzLvcxRrUGDAba0UFi4ZWNyqbQBjg/D41kYSpqanbdFxrPS3sQfe
gq2eq0Bfve6wcD1muWTyF0oWHlZfNSZaH7aHnzz7qt6QVkudxYv2+cBjIQAe6Ya7
cD5oT+9bJ4AVyxFimwhMLKifw4W7dEDQMvL8oREq6dfLYqCr8FNxMHdYwMTjjysX
ai3k4Tt69XPAv7DDZmqSe+WWNWU05EIumCIPnzUUzEZBTmCa7ochePFjnDsgd+f4
fQFCpvRKIiWORednbgfNIKdQnuAkq4h5kx+iHMQLexv82l5mE2B70C30ZJTzlqiy
6plKVx0GXbpknSTFQLv++VaHYvnqW5C3DfJzgcQIWUdcRmc7G0XsXs5xloKpOJrc
ZfkgfUZ5Tdl4oOSYyk2lr2Cds1obMz3kIYKTiM67liAxfLvv9IhccVNzlRZNihBn
DcyBgVUXtbJRUI2hirY9hdYTZgwKdH1AnHOLa+/xXJeDkBNdFmpvvESkvAs6NkVW
xHGxkERmkJ8l2y7cy0IQdytIdLtOzHC8e9cDuvB09ZTUYNXOoire4pupFFOF1gjG
eN+fPtDPaqhQBFOf+iMTYVu2eU49yf53ksQGgCABFb/IyKDd6cp8y0lEdtQlgKcK
M5nZeo5p//Y6qkswjwLV/WspcqSUS16Guvyivp42b2OaK9BJgqKehPQ8HmBgnkyu
YBAfMn5NDORc+KTxvYdyYehDnj0yrQ2ncOoAsZu9XnVJ7hJicfOgAMR/F8LkJMnd
UQxEi3VSIW4kYdWn2lnJ9wtXsPII0yZYKUUnv6biOXyKRO1C031Er5R2kwHgxCHd
eBzE3JpXCJhTrcuFY6KB4qzzizYvMvb8BTGimCxcw/hUgr+ZhSDW3IfMaaNij7Ln
xnmgr8RYo+BtGxfeVhVNftbP/RFa1NUsNLetlDbSmNXfYdAm+555biWI+zAMYA4C
YW56WOd3hz7AqWhekpLIVTBjn76IzlKY/c5RM6IYRjBRNUcs7hOuFjjSM5uX3OQn
+W7OkM7Y99VWWdFcmwkZ+da+uxjtDa8ZJwUmM2MBT3EDzHjOq3vUa5z9muFJ1Q21
RX8MDydGzzSG2PqN355JWXe82xCM6k53s5hieyA2e8Iaz3nih6UYVt0HryXMXGjI
x2xRKR1VZFaZZAUKjDYXBemL7RxpoFT3/RdAz89Ur5uoG897XXRRiUdH0vuXn4qi
06wkp+jzuMCSfB+59+0a+HbLbIRvaGXA24ZTpVMJX9zZOEK7UP2l8BdzwCOhY15e
t3MJP0ojtNijVyZHszDUKLpt1JaGp7QmNwTyhqREZEWGJYmzowCDe0NfhuAjfjSZ
iOQbYJ65/zvZzWD35fi/QZ9qk1viX4088JlWo/q+DwM/2qjyOLbsHWSI2x/9GYzi
p5t7jZA6wTpg1NqK7RYAV6RShP9kvlmiXaqFxn6nykX58ZC3uOF1HRxxq0tNmEkp
Gnv90mQ5txnQne47LUP7F/FRmpM1hfVFaTBVQmvBO0MQI00bEdkG/U410zl/SZai
+fKqfF8jscJ2CD8mGLGeb2B8zlYBD7ZmE7tYV51p9JCpMAXBcKFd3vpGxEE+BtR3
dWz7RuZyO/VjQWOO9wouQnyCJSeoV3u8o6wNe2PPfhbl060GJBRRlmwa+fJimq0P
3qt3add2oQHBk920Bogk3iGg00T9oLc/U9ebBl0YEPM7SJn83QWFjiuIt6Eu1eBf
B2V/bq/sk5GhshS1jHdVI7m8u/1zH0pmZtWsUi0UsXXVGHetANQV5ojQTMMnUGzA
SqR/E/+irZfLLoPWLBJiFB6H8PWzevCQzhFCqXHLLNsLaAIalXUzGppNtfGHu6Ar
pPYUKX/ONCWGupMONGe8WzWIjLSTi5EiK0GIo+PPyXLfiH6/T6qjV++c2p3JC94N
xe29hp6LcNeZHMcoz7iw2h4o2MYo7Jqsc0cm2g0UbrpTQcH3NaUz93ZTucF5Q8b1
HGPkljwyIgEHzSgCIiJi6l6r7z+08/RF1b/X/56BJZ6APeZhLMf1pyIsV7fOZ4+l
OuDtQQR1BwIfx4YOQOxI9GN5hxF5JT4W10SRdIFH03jR8Lp/2Rtwvod90yYz5gMz
hpDYPXKwjatnDhkDlkuSja2L9wGWga3gM9sa+EzImkABKVU0W9br3jEYxcu1lfmZ
UK6cidi7LTB0JC0Ve2TfsQNZFc/aQVEPra/o5i0e4dgGEM+FwHZIeUkgKLgXl6vN
pEK0qNrmGkcoh9nyBzNNb9uKy3KzWUUfpjo7qKJidoBYoqo+MnM2AI8e4X4SfYOG
M6gKX1uiLhSxsQ72wzSX9owSL5OfQJ2UU9LWP7XsBFy+Wwh2GjkJlOlfTJLML3OA
KG9uvZdJRY/W9wVUZY4WhK/aPEhM3VCajhjmDjGeyhBeLKcn32kovGu9gW7AO3H8
+6vqp/ZGpAfDBX4X05HoWrCLRLwH36g2CmMpFZqMGU2Zt8w6grXYFFsbYcVGLt4g
W2QmKyaGlWlFLhCz/15NfMoIAOIiKCX9GGfSoBRY8VC6324+j9l8ctteTzDpU+XC
LneGcxymTkd7oimQ0OXsnZ8fkYQKtp6IRARtpnjesJAnr0g7o7Iz3pyWDhjlrT55
pA5qep/jqLjtcd2Km1TIr/EfLjIVcKcj9io9pwvLNSEggKsr3aG7hGiArVE6asXm
QJffIu+0ohB/+oF2QRsLDjNAwNTtEJLsGr1oaOKL85QsZtKuOLIgMKue3Sh138ui
+YRD+Qda1LiXzYPlgix5hYimr06bAo+6VBpJy70vVojzHe+hDfLw5uUfpYfMUjee
dt6IzVNTkD0tQolFB48N3IPp1sxringeztJkEBgbUGYCrPf+yyA/eJxJpLBKvg+y
P2DysiDZiLLq/1cWmhZkdN9WwFY0fjCYuZaRCvckvYjjGCGMzRwqqsyKZAxrw4dq
o8MlbDgLF/GxyKV1rv1/AyJNxkAR1C2rk3hsMh5/mCif3hFpkct02eHsVIQhWJ24
ixXIu3wnTFFqpGUY34WFacoYyK0t8OcELjG6G25yUbOwI7bvWiemau5vGLSza4U8
8y1+p186nzPgRbrr7rgf+N1WA0+3BbVeEuzRGaPacaYtJZ+na8coYkHiGrEBdUUV
7wowrRpc9GYNYEJiz6p9fPzQdwgjbMQ+dJNjUHuAw8BJDgkNNNa2pxEUBYYqjGjS
Oi9xKNXR13Qyb0Mj1UqVIxbmzKyH4R5QfTgg+XJ4uWgc8zygHLZOzn8K9JM3yz6/
TymjJ0KdHl/rQF8jNxkrmhcZUoMseIk3tf4Q9NM/r/qspmWtkzYkbH+PTOdFR7XQ
KsMt1Iv8IkEpjl3rG892yUXf5NjNtyS0MjxrSgB+bnTEm/OBLckQTB3Uz2FkccqE
HSl+eZXyZ7XYxgsal0POimGLyNXuQr2bQWka6jFDqaHCfNaQWLY13iJjE1BzQ33s
MA8oZ9jbVkcV9/FPbx2iWCziJzuW8moc/w5iVXZbNFEulRIkHhxcApv466j09uSn
m5dryZSBBkcOgLANr5XMXkSwrBpRofCG2FpjEaX14i36U+mj7+OT2FaAPyTcXJ7K
Zq738kmJkfzc3z1HpEIAEqsh/i1DPsQjRgoiWr8DtvNGhmRdfn9+S9/gIgiw5Fsf
1pmQaHcPvyft6wjfEDRbd/AuSTSlH/L3FNg31XquEo4ZOMX/f0HM/nMqZmHTZJqV
E3dfL1KPcAm2N8868gMGKZv1nZYBGH4plFYaVIy5fi1b5wcq/xOIU1FUX258G3zR
Uhk2pVLZdh/4dT6QKEX2rvEU6uy81STfc+9DAMGNy5BHG3PI/LV9CE48vF9GKMFF
gQIJFsHd9aLVpklGhlLf9FrDGWNVzk2JP1tq09BG5tP58CltfZ5M3IZW8iQ3SjQ7
p+PfzczGCGmu8QBRUEFNOesDa9+VMDQXmEGGkASNHUVNU00jMxhMGRT5v0hIWJa0
7pmUUIbDJD6sKJlrM9Wezh68yv6LIiH1MnM2XPea0i0PO2fJQd/YTCK/D5rOLUMk
mLDUNjrqoXQGE0DYNsApSHHU2oSgGMF/mgeFnlrvl58Vtug8PTsswnRys3FgRRPc
wpzsolCnnWPpDiW35XwzcVXLqHGMC3lJWmoD7+NmLjQI+hUobAWKFyEOzppOSyR1
FjxFVC6xk2dZjDUu//HqUC86nOCpgdVbEQ8Ak1WHOpihC+SD1+phVHCYyCAhCVAB
Fy2ZRDFtG8S/P4ygpbsX7cORsXw5nF/lD6ZNJ6O9RgguQAzEr1uuZ7QQJf+AyND5
bt7r8xdhPBMI6wimr6q6y90HwYuQ1/7JO/7i/G3U1lPEmaQ+e2bv0UvEDAcpA/zE
yzy/HVpRI0P7zu39EZ+b/WASmG90FvaCdpmDKMqiexhGixgR/dMzyAmUd/CnKJYr
XK4pXCzPcE4fLRF/QT0/WpwruXhRnbHXVxPtiP3P7+Jpjzue5xxZL1ZlEFU28jUw
CnIt/ifk20xTHuGhUONEjZhFTOJgw8ssBivBObQYH0T+uMI+oWuFyeLGn+vMgQHE
PO/UCa6vwU9JyIY8TtzHlYH0MPsmdrjRQoZr8a+YRhwGiI7lDErSCPCGhPfC5ynp
wizZvAlBioCJVuC5YFozkrXt7HAvV7FwwRYyF45CGufdB37MFyTeIZeBU5GSm1k3
QEVjLUudEU0cKYNeStWLm/7k0B+KqKxtnpwxAxFXgINm+oLceoKxsTnLQ+v0iSVe
JDu9/Zmg3EUboxl9o4Hi/CKdMGhCZWwVdIF6pQTH63iXY35ENmN+T8zA7VR8hdcd
ELclgWo2/oJ8g5ueSrIO6Eb6AJeiIVkkvSMDeyN2umTTY2hfuIjfmNIvDPM7qwv5
mvk9Q63lbdTpCGjrRhzRMTNTEeW5Hcyb0Et3kiLkjkpFzy1nMWWbwYMo8J2dO4Vi
mIg85lvZXbXIpMAZWDtiP+aBNk3im+hsSJV5dZLvXtzvG62rHvQF2q7DYtps/XQm
GGMLopApy47OtxfjqGI8wbYstdQfRSfJEX52x54aro4bajsPcm2DIAF/q3pBWqTz
EzKhPr+z7YwHa7SaaYQNmg6PmSbcSuJLQTv0MRvCt7eFtS2teY3ALmogQuyIMEPG
3krnrzGfb4+4WUsB8T42Zi0RZoaFlpZn/OC2vqd718pCSjV4V9doYYc6m7y7AOZO
+ThiKAuwRHcp+iok5IjJW5/d1+2k2LIpTlYZmpoqcaRcVcp8o908aDwUJULyiaJ4
eKq9wMqAMDGV4pO26gFRgseMTp06P5g4nst38yE9Oy3kNf7kABbky8ToNMXYV+Cs
fhfNLBiGnpTU+ra2HmhS+Ln8yqG3gxlKQgdRI7lSO1a5TKc6uFD9TvYMVBoE9Xhr
z27DgF/UMZi2KVhaFoiRJwy+Fl9BAbwsDJB6AwgiUTSdFP/4PDbOK3VWSv2+4fCI
jGM/CnTbOJ0QfWRnHBRCFATMf2YQeTmAAwyFAHcEQESsxh3v79Dyu8p21VqLmNUJ
TZFM76UTkR0ax8QVoEJ6zPcdH7ZcvkOd7s1u2yfvsKhP68bnS2mvyBbXpBiPRnTU
zMNcEEhKFAdO8xRo4tmLtm+ZcbNez4/TxL1ZObtOQ6Rmmw3lraXvKErnONvk3SDB
zvduUm9+RQqnmL49ppBREdHyRMdhqBy59OdFoN9sGEDoUhc9R/u/1Jww6+Bfz5yQ
0s7a7MPZWoHqQrIVcvaqhJFY0e0tBUzgRbPy9kszdAS7pMkUoIwG3egTi/NkjMdt
rGAZRzPKIKniWYtfFq8TAJZ816RXsdpjz6nKedQXnrvkQ7IA/XB6/lS4tvGjEVIz
/hkVvdPLjgATSzOyTDNRzVZ93QwEAcSEFDnJGWsCySLL9NxHHHeBovco+BbPVl7h
64g3allesIwb6YAqV/Cf01bc4Cy8vtoXTHwrJj9PrMdpBIxLDfgFZ/M+ZHdho5VK
GYcraSHJiM0VZ8rZvR6TzazrTb47ZOJqgRGGhEooWeol9P61Y0IxN/80j8Ryk242
Sl++BCLfIucQbfBDhzn79u3mpHU/k09EeD8u9558ZT9Y9QKYBa6na+TCFVaqd/fD
s1NQzCumFC8ASWoRtKmeXo5sHt2YdyMn63DQPqydnWrE2DlzpOwrOaEYnO5pveqk
H0KyR1I7VJxfDV/wd/l9RyBVsuAO8ldz3gCvdn3NOGL8/ogm6tENUQXtEgCKnbnY
JUP/3Uk0zmOUq5HB7mi/t+9E32eVzqNT/zYR3uWl7Z4i+XpoSDuMH/ou8yGOJmhU
4FkJrZEikpqa1SdIWBY2aRUBOQQxco70xpak01Nm2pVFkPDlzL7boWKmY0ZsnH8j
TACnEmVjfXbIsvoDfoVqK6hWD0UDy+ssURoFRLPAslltz1GVuhS6c6OoTx1WmO14
Ypo9y9NExB0mQH6G6s0AGEyZlkTJn+0HmyxGHazPPcqrCyCiOiTNIguB64GbNu+P
BysOVSXeFO7Ekx3j4GqfQKj4tVWQpge4l/OyAO9OvNzbazDuhfLWnC9l1OaAbc6r
GuVRnbF9WauNWqpIGLCt+KTdb2m0uCXnIXMsbIH6YBLk2t9xTHvhyVrU9HSes9FY
JAYS64xrmzPqWN+W2MNcTT86QqTgOzRUY49aYY21Q7kjwa83rP3ms3hpBl/0+MZ2
GrXWDlCcxezbyeX/gPSCFNKzCFyLWC/6hS76PIB8vDysQCD82Yw6tEjkIid3LFVu
dr84uJLPhsmAPwBQQOQ0UQA9aVKUSWMG+7DZ4paw6lZ/j9EJ0eGeL3HlPmHHP5Fq
LYgEuSSHVdMcFPUDmCNJc+kHOeZB7HS4jeQBmQv8ZX4rk0CDtmDHxVSTdnsmLrLO
xOtlZEfCeW35vbsEr6UgNmJcugshW2Dc/9FH3be14RfVk9+yD8I1exupCWqObCy0
2x+FIZFKX7Zs8IeG0IZdSN+tFLVcqxflFnepgcESgj96UbbZ0YH7QTFhfaq7n7Pf
bMaA7mfvB/58aDXRgs4DM02KHeH+OPSL7u5PXzSPy0KCu7gT5oo5V9IOt8UrdZtV
AhdPCYDY3A9iiY5/vzlSvsUQ8tnmNFX4XKV/XPAwpGU1EMLori12LlN1QOGh88fa
HykC/1De3D+gsMILH8KX5QSYJ/ZRSlNW8HGelCJB6wIBJ4ki+sk2uepN6puUJBUx
TNugySgwwmlkcGWiYjjorC4ziUKgwCZJ4OimlEXb2QXwB94n0y+mts9rojlXRREE
cuapuovVtPjqmnOFTNpYdth5TmV16CBPKSJjwJR8/duipswez1fizVO0dsLQUMJ4
px4je9/Wx3CnhcXwUsV41lW9W+ge0SvCTwrAHOA1JbcHLNspJcNxN6MrcAdI3Blt
l6sAtdDuUA1FsybJt31Nj8NnZEUBNyA4kzY7AEuqBzlzoRqdTIz9TodD6SW2LtLj
NvYpJBaMeTABlZVWw181r9/CWH5QlSWomJ1kWSL8oFuTcLjnyeKfyJoxhFOoakZt
eOZhKbHGqL7Wp2V/biWenCt2qV2ojf7gcbkea4LfYuln7+yJFCtBtPC+8SaUzF80
pjF3v6jRCGrzQBe567hSabCseZLVOtvand66pTWvvITvSz+nGGeHvNUOBp5mrqMm
98CtWnQ50K6Goo1UosxH/Xm8akCRe1J4TTFyernidFFKDlEuGn2xNchnJEL/iXJ3
JyYrZmwtiggDoQmBlWLmLg11hycjSwZ/ycUzEUe/CaMG0TsmaRL2T18DI/F35Vze
KgqzniCOY5fPm+r0tC4gmc6aERhAuIQdj8IXFje8zw70q1956osgNfSgOLfBwabG
BvfiMwsTsseqMYMcTqdhWsQFdPNO/XyxQ3aSTgvKOn/3tstJe+paQ7r1jIb9miPO
+hrEDGk18b6RJNGLrLArVlnWD2FV+cnn4cMyl6I6T6Cj7RFtAqjLzaJwEUh2jXRG
0fdA8anp/JdEx3G8JF7akkanhM3Oqk/Ga84TgoGKiAJiiikt33gc5TVmBg1A/Ov0
pibYRfeUmuDCTpluZrZq5W7hpsHa0Pj3sHr0l/bMD0Ya9wVVKxEZPlur22qLXYxF
4ydGngbMv0xhiHknhJ+pBrVyX4IQGNzT1fpand7M4hpnB6cyhgf7h1986REjfYUM
QcOJbRBIgiuFLUH13Nll4c0eEuXuSHxqsWuQ3mJXIhdzQn3NoMLnm5hI8SXMmhbt
SKhs8zdHR33ocbiVbhiB8UmygykjUFXrTpIfmdmOYGNGUszz0wpgEWJgZdvKzfBK
tKTmpOH+rkMA2bWuA5jaZJqHY/SGZ3+czvbMUBKDz2d6VfW6ATOcyepSlOkDU9j9
yzMOU4vFNAdAwzLhIhcptwqGd5L28CCy6cFnlJKl6GhzD4Iv4UW4B7/xvctFBf3g
ZEC9+3f706T3NU/RRoUfYdcxrRIKlq55BeRJo0ZFj9H8VbjYbQKWUJ/2fmuxxRTl
vsn+2bG7LpMcenxpQS6XbCaPIBI0aSk/v8IqwlXQAqhqTCKjD7IZHbzVNI8dq4bh
FBn4KMAWNrcpaBtPgpeIHJ6EY6TxRkVZPPByCqHssdMlC1IGNGJ//OHjnWWsC9ae
UdsLI06/XjEveJurCy1sVmTFRb4YKeOzzttIx5TfxSqV+G1Lu5YobUIYdKiwvATB
Zkq67/VjAhUFHMX+68tW3WYAwkSNzDaQz8Nug4WZda+Zj4l2F9MmmPHRmFVwVSg8
cNASHL53lPw2qg6FoUWUAWxObPSAdONh3RvONDLFCUcIIerQQ41Z6ZcuqIIrpo+w
IGEjkNiPbTahHTkzwDXk7pID8oFUaUOoqBsw+R7PFAZ3G/mZGPEY9L6DLhBUxe1q
LIbP3HZKN8Gw9ji0GYivu3PZD7ff2xLkfUD3+GWP+Au5vshZOeMy1EMaKQlOZzFM
VlUDJSXlsz60gmUonttCYmkxkSJaBwjOYcTUhir+fWCqmqOIDzq2nkqf82qvyXFQ
jeEN0tyHngD9D68sdJpJ8t+yd7N64WpoV2l141tdc+yZuhxTzkL26ghpy9SdqPfj
rT3zGsTsyVHO3eGJd8D4Ch/6gGaI3V8o5W7FuFypN8v0QRquhvXF1Ql3Sm1C3o6g
R0VNzwaEOwuWZMixHyhG06stxCpfYEY6o7+7LfVzbRJHLke1PsvMSpPipIwJEtEN
wauiUFCRJDQmYkC0CmzvT5TGniBmw/7+HtSvW5Cx09gTx7EW4k4EoZmQ1xBSmE9O
8rEkVYCjMocOqWrULkxlyMvOdhAC3nuzIZZEZqtMDy0h+BipocuBOhUbIvDXrAI1
Hl0OINTkZymgF9od4ZnAxwfQSqpCqlMvHF4ET6a/VPAkcWPBMf96i+x6cuBFFSyz
PSG1lS8oXdOqLIbaFvJE7LsqviFwPjvuyYulVz3Uh5W0ZtML+1GgO+6pKlYlwaY8
kHZmZFa3ZLAQrOTwOxNVDtLHaD8wBNPV3/TC7bqX9Pq3lO6sAXT5sOBXKvPPsiQl
NQKQn/TftWGTbUzvuhydsRUDReFTofIeJat1r6Rnn28vuReb9zwcslNBdvU1cWGz
rQpo528Uqg/tB7sxwqqNH6nbmwxYslMuzElP3uUdwhLiHVCIcSu7CLFi5TiHNCuz
fWhrE9EGbllP9tiOGoCnmEAx9PxMmqZauUncTUKqBzgBG2MELLWlcBBw46d096A6
+ZGvvxTtVSeF43Hi6dIxyf+J/nm+vzOfW/t2Wr7MNncz0zxTOfO0a1PRsKJGM2+X
hGM3gC508qZf8KH2QkZlKD/UFLomgQVMwO3+hOSzuNaKHUjLkGPHVlmWpOesqZpb
Dd3bO8YKUlBo+fvDfzhsIeexzGrhq318hlOJHh+f4umqKaCQwBZGQ05NMoK7FryB
u3qsasYtbemMrBmL5MrqKjFC9PMdQu7oat0JHWAMykvSa3dPX2wXReePjs0JuYe2
d1mHDyaHgOn1TKD/6uQ8e/+q0++Q37O8rcT3W8nZ1h6BDFqeBcLnY86NTlodXWcz
Zaip6QvixCPw/uFH6mk9wUOp58SPHzkNnnUvrGDj+Mi/WB4Z7PxPpWOAMWl/Qs+/
lBQ0exeA4BuBpvjQfO1D4wbWJxf2XvNxCtcorAkUsyBeRA6Naz2xZlhz9kO2sJ8+
w0UM7u+HIdEgCObr1HIbBWCmMn7kjyxQsBqqr5d2Xn7WUsIxbFdZEDJZcEiC2oiG
uvbYDzWGnJWPFEm8xN+wajhqWXeX6xooyFdaBhEFQUEmm5BlmjeqexkEDVKS2Rjo
LvmvI9CNunOfYj/P6ou6pay5BrCKerqN8/dPHEG4DTV/ahppprcXOhO88Q4ku7SC
dLS1gSTsRK3O7+RooPdKmFqRhdqdL9AGtuaN1rmlKO6SaoJgZe0BpWD1coYTimxf
2acJ920YeckGpxiBXtxtxPDO6S2/3sLsvPF38tqAlTUaaNPxA2VIomb+YHuWUswG
tbULQi9NwYgHrDpHpNTfbYdE/Cxkz6Z9SZQtA/sG/yknx3bRpNZj49TN3YAw4vJu
ik2E4BnLQzStO2oKBP9E7qa/Es/tTR9ED0mgRsbuz3cqgQJzFbJDxhLaOdzgm6V4
/zR1ojIV0iGBBqSNSHhoR89Cx13RYA/137cZpErQP+xgj+uxl5nJxeBPTFPXjwku
1ShYlFkc1vAtwMcch6nF+1X8l6bb6UPMqSPSodHlbB6psKi5X+wkjQ22vTOy2Eji
EIu1clYuGJU2s4zNsNcEgkFM2oaC79qJvfovjmdbLa2E8PrMII0PwTamwToOVACl
Om8VtSflkDvKeqNGBtwzacjUOnr+kIR2J17y3jPmgSHvR2GA40FGAkrhorIbNnXU
QFEXaw+yDwoHA+NYX95OTUC5thix3KZikgNKBGeC7XUvq+sp6m4LyLZP6dsfyAxC
W8HwQFNcWwmTwOqc6wWaplynpNSdFy0fEHwpNb2lt9JjTDg+LjE6f79K/GXKKmbK
uOuVABjPn37Vp3wkGo8UI5WwJ/DM/EwAOyAArmZTpQGUhw+/IbsL8d0/owlcrWO3
ZYdIzTH6tOQ1/14qyBMb8Qjjp95RmEQG3Aou9TiscfT5746+lMrxavkPAzF2cSxS
df6NquGu9zurOVh4lzLzRWKd0G8V/6TCeWjnnkni9NE9lRaCrdnCPWZQb7qfpUZT
Imv3YnDaYMNvD4BgNkhpd/LbjpK7R29s/vDR3UZlMCHAY3bqxSglsCVIBHOMfv5I
bLkL5qWXzTipVcpQIpnaps5KI1MPSAGVJmsFTA0NDrtEDtMxPrz6DMHPmHqvznce
yUWbwc8OpSdUzoeVRJVUuUEiGam/1ZLIhe/iNm9SKev4pUIysYWZ+KN1DHlm7dSN
PhFeGxvuilife/lIOfavJyaiQVq7x14xyXzvkomtMG0NUsKzmzaVj+e3yJ2T6UM/
hlSCujfoMApS49puAuVfga4a3lBM43H9HiyJ1Y5hbhPaBTftJPPqFBdSugA8uZnW
B+agFLnDYeGDRTX8Bs0SodQS0/2sfAPC0Xy6nDBHxxUHh5N3ogxVChulXVf39ONl
L14eyaE60kY8aEogUmvr4rCgoY180gMitlDRoyzZzhLj2d1go7Y2HpWJZyVEZzQN
SvR55l0ifGuP3ilV1hKsXF4CAIl5SJVheG/UDjU3WYwCiE1dcUpVC8j0U17JxWJl
oVv5kA4BkQv4CE89hO+k1h2oZwTwCjJ6+vOBisEnEVMp7PmN71g517Cfakh08JYK
Lfz4Sd6oZ85ofECDVULIazGBPePyeQh70l1Lb59dGuGX7OOFTw/6ZUXpiJXi2a80
wv3Q3Uy9W2D8l9JPBpe07KVT/Fx+g6LcD/O6rneVl1VIDEscSeIpAcqgQNh8HNnn
VODQcAfotCAeEfUH5/g+I9qg0U04lyJES3OnfioXgvBPGE30UlAMKLX1T6v4RAfL
wjBAoXkuuCw/TDqfyb3ra8hl/5ppqhFWahBypWMmzysgWRlHc71MGCy46GaLLcos
Vg+pcjZ50bpbX7RV/LjK+L/wc2fOt/+1P0O4s+O/iiTVpLmYnhbMLMgl7fcpOtny
qu2jxFFVP0SGJJBR7slxwwYVKORPuJvrdBmhLTL55LqP+zOEkiu0y0gvcb5Yo4Ym
SlCgXVz7f5yvLIgOQmUUMa/0CzdfUQNpobABimTUrD1YUAxpN958cjtmxRkDZvLw
6BxNIAp6Ypl1xe0yePYzRpNwhjOCzHIAtmdhCyQkfS0VHfT7jbNttrVgETExv/Jz
UvrYCAOtFn8SNMaAbz+R+dZzCbTF50dVAyFnwrZ8ToTmTbk9hx9nf0a5szPyFNOq
DX/LvY69PneJBtdPD9uMih3q7BeS3UUMTzvPNIXW3TXnPicVHOpvuL6o/5Q2YUTk
EypksNmH03FI9yClMpWQlOS40JgxStIBYXHkHwmE2133TawmfwKhoPQOK0q250sU
e3dhGKdUqZuVVJL0Hsclzlux379o/FcX6A3BH7LzrFhI8tgbZ56y2FkXq1reAdEW
GuyzfX8mqQKDeXGSKtv5hgTCKJGL7VcO7jr5kSEeLpILelNsTbJMMo/PuJVcO3sN
xV7E9bkF9aoRnrtp/G0GI7DM0RWYMB0xUtaj0qNro4nHCGlEkWPgoBkLWcFPcG9N
/ItXi5SQO591TXAv7mBVWAr2TOLz319XDPDJ4eM1bFBwhi8sJnvOxRFaBXrB3IqL
fDVzN5F8FJDIXkCDOnqAivMTgBaFYXDpH0Rh8Xii/ATNrFRfNyDp+GLsmblMx6ic
qzkzHk5iadh/l+6x9tOVJu+QG7luUo0zsUeCWOU8VRe06gnrKMMRdreUOJPMkf/K
xp/l26aiV2evMdkI6xBsg2RkkizEzwzCIZsrpix1CY4BFMUFyOhlW8Nl3IWd8qAy
LG6sUA6qMrvObKbINHrpukFK1zsukFKLuc9Sxd1Wpcw6CZch9QrC8aV2ktS+DjNP
bivrLZOwKQ6L0tJJoPxyFiHLLjz/3/GVQQfBeYQe/rUeHTp4LTYHQLURy2J1jXiR
ItB92+Yo4nt7rQC1tpFlmMYbEOY8uobtn+x83Lg9bqa1kmobzKhxXWI2iOT/3PgT
YKFTE2plMGASDeNzMIP3BHO1yWow9omRhwmfev0we8Vnf2lESJrO1IRk8qrvfIIa
0fvMESUGGLP8ZuKCkKgJN2pEr8LROlRb9+01hgQRMnisKE5Hfk0zXoAB6FhQlOBy
uuQQr8gFjAgVaGw2QnkT3jWzN61zWNyOG3SMokfQesGTRisIzwhNnHRJJftr1G2A
3ajMMF9FuLK1JWK3NIawU/SSa8L8IYLGyLVR9NzYsRp/hVw+gZpQqiApoqdylFox
/iAI/iA2NVtVF5IuFpxy24zezOtOzEVVLJJO4xQ8A/GUmxvHM95M3tV1AbeH6AhQ
peMZ2rR9QSRZ0ML0jh+jm8RaMwXYdhJImTy4RV40j8p3UJR7+xt2EmjcFa6Ucv60
B8Pbv7jhNM7/6QHNwBqu5OmsFOteIogRIH23I5Hvig6PAerHKDPVyg667NVRujJK
pv51UXnRmwrT4v70yIzoYUOoIu07KJ2XwbJNyfyL+3LQCnvmXvb7kiNWDB76NOHM
PdLcnLR8hYehROctU13SiSd9EGwhaYsU/zKpc/SCAFHXssrKUxbWKirp5uoqnBiN
m7/q6wyJglndyC+yLWR6F+vSLWueX9JrdlCAGGxeIKMHOlE4ZLdMpT55Hl6Pw6BU
WPMU4RV5VsinZfcBbIQkj5wc95C1+ZkqYM7MrDs8fkgzBXvjp3R9nfvgxBmgY73L
/emy68HpcTnaKlVuY7ITQq7fyKvVRwPCTlZZT4rSiuiISL+2yX10HNx4gc2G6AHU
WWYxaR0D2yCQB1CD8asdqI5IqK5TPh69dI2HCz6zPH8bd6ASDjh/0Sztg6s+U0ig
mWe/7f0ZpbzXprjiHivUqDuIbhyo6Mus/1bdTyRWPMvvNOaAjQ1lLoKpL8GvQA4S
ZsKlEMZcbM8HEJ6ey3UeeMXti6YhL2d/Cl0xgAZku2zTPQ1+xQnQDeR6IWs1xaCA
Q1/pItP1uLhQwX1hNPyY2FjAcv1SpPDURWFzKwSU3mHKzqxgDEqaquiHXJd4j/Bp
HCHK5M+iwOGZs8fTeaxqs+fWHwTdl6v33Evhue6N/WTy1MDOeRzjzNtw4seBtbuk
XuT1Mn6t11fnmFvKZMjb4O6o4ieCI7R6AbwZOLuZ2SjOa9fMLrFh5jVuJUPR8J5X
Gri0H1rbpylriHawCSux9Wh1z0wOwTk2vE3mtK0Xqk1jvLONa+aeqRoULGflGmYV
TyFNafLj+Q0WHqAFW7KY1br+8AZbCp41PUCL/IcsANTbnNidwTDV1BN8th5i4m12
2m4SGCpfjCtlz/h86GVNaAipJYKhPKibRt4YApIKM+2Thb6wzAG88fID/QO2Crhe
RTalFZkQ3S8ulOgX7s0D2y/oTaH5pcSvXgZdyX7STl//C+byv9x7M4/lFcG9zPvP
ek/ZcY6YKrwh0Atp2XcxFgrwXAw4hdwnBZRIGh9CX0vUxugggckLmp9xlBbqcFAW
NQgNWSVMQK+N/9YdKo+HAtF1zXsNNez4aEtrF0eJivGFslvFC3/5hhpsghZTvydL
HwbyjivBoSgXkzPG60nm9RITDVx29Q3z9VONbm7Ygks91pqqzfJ2NnA3CN1iTlnp
G+BSViOByxjADBSiyohcdtxMpc5ffjjADQCw24/ymxwu8kCFUXWae/Be99DrUumD
G093Iq6Djx9Uf5R3+LiuxutdC/9m9uho9J/Nt65GX2ZsmTRZCmXw0C2TciZM1x20
LVjwXEnaNz+g5y3aMuVlrHb12tc5WJjtQj8ofWeLUQAMZhjCqbgwMRIdGtoCfJ90
QwBoR9UShnwsv48n/mmj/NEbrqLKye7qCbJGcKlJTK3WMS+/VMfIvDc/HZDjSLmG
2PBplIQyRgHq3FPhJ88laTnRozh5vTIBkd/8KepI0yWvp+F4gWPOxkLcCI3MhiVX
aiAfHdfQc+XyDPOcnzN20G2+k/HEBPcyvlCDDf+2YXXoE461O/ndI1K5N1Iq1LQ1
xVObw5VvCRevilyF6nWA7VUYs0W0SSuwFqwe55A7yGzRtDsvVVApBMTH2Qx3pP7e
HH9Zcrx4yy/0CZzuE+PTVIfe6e0m72RFm6aB2IPLy3hsiaYeiqzuKkd+FhkmzadM
ugtZiz1QDU0NtcexM4ujUWuMqH6XK3JzdxCSu+n/eQK9/nJlUFo4gGZgfIUNy5Wq
44PXKxmfcJgDIcmVi5f6xprWCkbM4RtNDGSuSglqMdGtGustAYQVVTUO6Kc2yObP
CE5w+olG3xSgOZdY7earWHxqN1a8+zGUqab3tMmle+s4FusPu2wxUNBkw3TjgWSc
0gYT9IWRZYrY3HxMMu6PVqEWZdulHDYiH69IKtu77k89biiWmfoqKL0oCkLoBbao
XA0zTb2K4Qkmdiu974ufGJqzt3/7MVbCGPXH9X1XBzClsPYQmfNWGJ4z/ImOygZD
+Oy7Q8oV6kel67UECJYMpWSgz9r1/1tgzvzj0GDr8XK6kWohKdZVOYSkVnuNkSOU
QLvayMvdYJiMU5NTToDXiwz4eUGlSra5AqEItmBebs2UnNeSJt7uCtoDO9du0KV9
FmrNh8n/p7ZyrSbAmAGbOLu8uKkS/OwKoQHNwwiSGDkQWAV7px+kBr9BIIXHCb0p
xXkJ3AHOzYNcv3kwsG5pcpm/qBwmIAIRJbPRjm1ZhBN7wOEDEG0SoifWjejC1Y97
1pEIcVP/U243z7P3QjhROJMDr8MMG3IEKe61tpE48fPTw2qbsxI/fbjorppnaosL
oAneGd/ZeG7H9whejKqQp1dqyDuM7qbKS6BuaIyL8wScOn+eDXVNGEipbkvcFSup
Oa3Ty0N0bH9fMlAu9CDPASpviwHTO3t6T7nEvQdJI3bz2SE62e6GH1tY8+jeB/g2
SrFqhV2KUbfZB+p/1G3QOjgdEQiOQ8yTPXfnFn8o3uUygrF3WU/jkD3Dd5Il4H8I
zI64p+GpX+gc8yskAc1nUu2UzQVKaQVuX9DPn5SxB3owuzL9P2/jaNqqvxTIzmw0
0ty/FQjWzLaZGwF8Q9p/U/9m+aCqg2u1wl23FAOBlUeT6Tvv0hcUO/zdqwtCWdUJ
qbC0CIN+GQ98pcgXL41/mNfTRLdwTkUEr6J9gNOdZlOWeV7r+B9NwKqyk6yd+k21
pavQ96wpDaUBxp1CZs+hRhPN2R4556LrTxDIuA1w3FRIhZr1QyOnpXI6Dh6lrw1V
uXlmgkQKF6psY01d+G7aozZPIS1+nlPaJzoE0nu/HmYMnTAvMzIZW0dtAaihmTv9
TxdJrmFbvWl1WEAnGDHCrnLLxBSqKfO0E9yKHMoRZA82JuqnL7fpy9uQXHtwoxPt
mMABE5YBS4nmQkcwl8pdUbxGxGHcXTMF+pG3QKiWPjeCuK/sDCaxQbArIOoFMSwQ
r+N64/vJCIeO/JT96KvHjy413VYB/HybPVZRoI935iBV+UaW5xiNZg4XC5sJJCFa
Ioxfafsx2/ewppnKhVzbrob76JPZGvByrPF/MEBaisw/Casdch2+7DgVUNdmTclp
4WEk4pUuK+FVuGRXP8BUuJI0NRiiFAH+aa13jbmo3XLBAWFmtdu2xjExxFWVC4fj
yY+2hiRAkRT3FkobiL9RV2qMooui5oYY/6ftlEcmXCKqdChQBkW2rQUXgdHiXElO
Yz1Si93PEaGy2NPXGvJKVnEuUpRGSJx8mgZwHuZwq7n+0PAwnzKcTqdt70AelAJ8
sdWFrOnm2mw201e0LuucLtl9PDd5KPUHc+I2BFsKCWkbtSiZG69pQI9INNys/cci
tqNGJ++yYx9tQBIyK7NUmTRKRL8VwLF+pvJD5WS9odHTF705qENehvU3TfZBcudz
vQh3UODxRvbUgOxBSH507UTLMCGybw2x4tLdC1V5plabMvNXRb1Up6qjATcWj1OL
ecehSrpYKi45cUvSEHTwpR8U1o66DRJ7487TZXuD8S1UAN0N7i9Ay46JpH3QaecO
Y+bOa6a3nbKUhiBL3d+IhFbuYTYlvYPctix4PRTvWvTv17j9P+sQ2m3vndMt/B6b
3CdSyqR4FRIS7EeccLX0WP8K72ElH7ei2j20N8cfstATcGH5aw+xQaQDri62B2vn
JXY5fmu+DZYvztBGTL7eXAdsrJP1lZOcOYKHAB+matxgJlsSLveDMN7jJU6ojTkL
/Z6zCGyaBDdrCCmlENNq+755HBdQM2Y6sgUQv0tVFOdp0nTC99iv1sUW+30ipNsB
rHqpRk+fPC4yONt2MiO3kwcY3dFwmaXABc+6fGEu7MZ9wCl5qcUSNziFIQeIXQbL
eGJMCDwAm+Go/wWj5dGlA3qVcXuZcMM5MSqFiQrv2JC25FE8W1Skyzbd/vP4lOjb
JiLE2Yz/OswcyY8IPQ8kmpK1hl1O0uMu+vkKfsb5JPZOlYsUoSf7b2nzcAtLtEtX
EtxyhwY+XzYOJtdd3sxYEQelmvPradCv1SAph/1hVKI2kK9zxK6iptsqqMeidupU
/C/nuMW+yCRPO2q8OBbxM2SW7nXS8LfLwWD3e64wQHkETPGKTTMP3/eGU+3bAXx2
C6urhhqKTazN1VslrXJPUDNjDGZFkSb+8lr1rw+C0z2Oyp5pwb0oMKoUP2JhiBSH
1qvTzL6EoO8cztrHFBzpsCeI+5YsgpHVANtP5R2euOaLjt64fzjVxkU9sBpIjJxD
2gIIoJk8jp9KzAE20ZKLTJyQ1sQGicpAqmh2aJhvG2VTBmlxzaEzeIUumIiUVU/x
GWe/IphSv1O8JjQe+rPgdR5Mso5gScib9bEHVl0UY30qaxDHaoWBlznk/CHGHGI+
RIlt6lCKYTuPSoZhbKiKpOIReCkscdfkt2aEJqNquw8bmkqOO560KlHcA2iD71Kw
wAPwGbhb0gPGGFDuAeztBlI8dVLEqH3gnk1gp7qq/qFCtdZYMDB6uv+q5bz9vMWS
zcrx/pQF7+k6dt0nhtlcrHXivXVJEb3bHxF5JCHUqN0ySK6OxLW6+3vpjpb0EDm9
Q8DjAaBKEvA9wIHcD/SMNCS7b2gXy25r/gWdSMI8w95g9rMo1XHdSXzEY/5k0hgb
Oz/1RgQoQtM+uX3KvbqQ/8BgLGKFF0gU6fHatozsyaJr+SdAGajREUl/Sw++0dZM
jgvj/+JQk9x70ob06MeeRFl472epGYv1+K183Ib78SN9iSNb8y7v5GrH1pgYK3Td
uxxVbKF7oT33xSDty2TN7Oul7wxhKfLQTINqXjRajBRnEgv2iaTWkhxCplcL/Z66
qCfBJz8wfFYpAjbRMT0PGljXUNRV05TzGvl+Y8o5gs0ZTjSOxWaZ/rBko9vxi8ai
QWao4aEeHmpej1RYo8pIO3Dlnq7J5Q9jx7FdcHLPUb05h9J3HkJ/7haB4axwbrIy
vp/v0DR6GtKnPI34Ns5f5hQZf4Lvo/Qoh24LAx8xI0gYKcPCynV4n8oU0rYjz5ni
aleR1Y5QfaAJ5EW4O71wkW7XNMsLpdQW2ZdD5HsPKd43uXG0kvibKGe49zSFIDf2
i5J6Cnaf7U0UHcS8zXEna+9lm9q2m4SPjXq9r2Iz3qFboBlCkR0VQ7Q8hs9lwaLQ
uWlBB8gIOggdvWwEfoHrg3sty2XLJQyPVWFPophxHk7JEHBzlpDB6GdeUbGStNAH
lAQePZqCW9lI4I50bV0+QgdFRGGLKXvJsIZ0iYoM7XtsNab+vNhznQFOHcmiUweD
lPPsx7qA4PxS/gNufFRFLbCRtQDTS/AiZzUUmAAAisxSryuu3HPxGfsuAtfF7rl/
17QuVpYN/fpHz4JNPAY0AzIPo1cHfswv2ojlQIbXes7TpZnJOC3QUrrCGtSqFVid
yrR1uNRBByDTEhnYQM8fzWADyUaiUF456a7t7ESbdLunNwgqxlyG7AmkdkLE+JmJ
ZSIDTRlcKTE2qABOBxezUOQPEIcKWj0o9XaJbanq4OJLVbvB+A+oPSHHTVXuFi7d
i78iMBzVoD+RZuyXLQmYk3y8UCDkOurLAGmKDoRYZZvuHvkP6xhyzAzpDmkN4lAH
rZRVLjpPN8SQq/+078BnbimYctW0uACKFzszPBj/gLwkUl+YCa+JUa9Oje1P9oF2
++4qNV32J3oXTQzkJLzbE5QsnecZ/C/fV4WSN3Kk1iDs/ZG8LV/aPJZNqywONzeV
jyfr3sy0MbgRWXVJQlWXuXO5Zcp9ovVVoTuXU2N3Rrv1WfjIBstPQSlIbctmFjBy
rGrtVmJPRQsZRdY+Ez4i7ZojubAfvbsMac6lNcbVPcgqsIiLT/S82IBDajM1fQs8
ctKEL0r1atuenSSz3jGGVD7MeG3ftKGQB6A+3WWnRDpCiIDRpnyup1mX8s+wQkNv
2EhHrfXkcSWUZjc8KlAcVYu2KHm3tdXAi746f0789jC6Z9MHbIQZV3RwmivlCLYX
Amr0BQT+Mhm/+fx3QG4jGZuh4CGRtoyDHK44Lcm2zE/RxXFkYWIbYPxJZgBUCCxK
nhDS5tyuO9gmT6zPylDKpFE0KFJA30uHK0hHR0CuI2fhBcENVKzJs+NFDHvcaRV/
5uCYlLSr6i97ChIxw/DIquCwn7GtTHlxhiZtftC48o0AWeb4TNh9UuL7VHy0UWge
QeEfW5MpqWQbNTXNzu0WG9KwPv81/IX7abSwwp8Jca2C7wTWwXHTk8BQNE1/pss3
ZUQx9kpD/WPSTPnyCyV2R+pYLlT9UuNdouC8NnT9sw8Ejik8kxWkBXvY1yytSWcp
7pk9EX7AB8cyNX3nZfVpg0fhth4gjTeuwMk1GO34QqynxebeWjtcPxpbAizj6Il3
t8IvaNG3hqolXf1D0RxUEbfs8F+3+lYHN7XJAtFxZG52nSsawG2n84kl91+bcRHZ
LCMAmpuygH9fEKZqNkFDc7dsi4PZQrabAosBmcmUEF1paUlbO6cBbAqJAcJ2UmwL
glLJEkqo2ifbuOauKPMm/WvIUd74aeOEe/tU3NaYGBm+eW6DTQUXkSFnurmIs9Ga
uNscrwXe6tiC2/H7x4NVoxggY47TRKyu2V2SenAdfKVFP1KFnJg2LqdZGZVjOrFg
R/T07mPm8XQS6xY0kJqymGJwXjMrs0Y5Um8q6UBi6rFJsj88zV8zXmOg2KNRjc/t
RSAp3pe0DLATsWcvxm5sb5CEqcqkYuOUABDsA8337MAyxU1Ewc1slRemcAsRN4NY
0QrygwI/esC6qCShXvT7xDcfbvnw8GB1eD7Y6IJwXqRcJcHFqYppD7bIsFLWFrU3
8dh/BkWe0JWB4bSU9wVMxeJnuBV35m/YBfVyB283BF3B6ZsTFYkVBI6ONcclzQoY
7H3e+lseKEuHxRB0IkHetz62PtTmjSXZCE6bzjaxp5GHMWUHWaRaOo43kghYwVbl
wbDmaXXzoQ9vwre1seqMbANySA6Xu0ChNeGGgJnZ7Wo8rExMPmDFer6jqfyXLLOT
8JvJIjqygnXa9WjZrCF4T7Qs4fWH9CR0pXze89o/d8UhJPbwTjjJYoL1R3NjNeTo
0cgrZnTRPKiz0FJ91vG7kEO+2EDbU2IysK+f5JKjJTZ33TJi4fKsV3N3Bcp9rEqv
uwDEMUyXh6W1GivMp/A0RLyjcNA/MYOkSQ+uF73oZSPyC2PNjs6BcWUQytpXcFBW
dJNSmSta9tGP631JCvexubTRA0Kqhur6+cxk4yNMI+HMh4/8J3iC9SuwAS66YxUh
7gyON9KIQITihpMturnm0L/PTi6QYmGDdaY79gOhH9qtqhC+SAGO7awjIN1yMn7R
Cv9oQLLx5eMqlkiuMMQ7VQI7tUykT0OWJrKi3H1yif+veQ9ryJ7Iq4Et+v1hQWoP
dsOWqjaZLLcinbqz213EXWpGhLtPx3CL7fcque9CDfXw0psWU9F7DR9NSX2PRLTK
g9AQoIwCw0bwZhFpmCwbQ92kP5LXCT+rSyBQUIEp6EJ8Do6Csy8QD8G3kFxUm5cT
CjcODKr9Rzm1fsPKJ4LehSJTlb7Vid7bF7V+ric//G4xhvNTJi8Z0r8ilO46zlGS
c1KBAM6lKDfLphLMtHgnUCsv5ZOiJrwHOMf90uh/d5h5u62IRZbbXM5/L9JjDM5L
8fGvbuOlx/akZWKF/Ju8wSsG3uSnMZ0JrR42qcdQxpRTIFnS7fQvlmXaOrg05Zsc
7INk1hds1RHVkWULP+s/+FmaWwsPIXSm1w7rIW8adnm1il8LewPZNiUqP9r4buvl
kaJZMbctUzwbh/XUqSIaHxnZ3zTinUF/43eGmtKhjZPyrbAEpurF59CJyixZzlNn
mNskK0DM3u3o3yTkDoeVnYbetjzRuUnMrVIlDBWtsjFbGay5DeQs16Inozf7+IKE
268NMgX+r/GM/MfrXnX6HGMHLPRS2RrPAhREIbHdO7KxrDIGXyQYW1ytmYoz+au4
I8zevnC+Q2rfYaDLKy8ydBd2jV9V8B1AXEW4WDgWtycZoMNAq43rerEOrNnLAS9r
6tbTJ3RC8gH/ffdvIUDVRPFC69xXk6dVTLxGjEeMRWHf1D/qoPuj6I78XTDhRRTA
Xb7xpPnREeczynsKDD+Qc0f9rcWW/JdY95tb6aB1WLxSq2/2WhUvvbwKIOSu0aJ+
Hy/oHoWu9Fj4EyPkMDBhm5lRUIYL1cvsptWTSfeh5Y64gxWjf1yJnThDr4Nz3sOS
a4ubpsSHiFQ0L08kRzqTyyT8BtDEIXfz2l/v7IiGulFdVrAHD9dYslg5i19buMZf
01GpM3bPi+ApKeqj6byycKdjkBr5l9ujMTAQ7a4HhChYmxhBLf268JOXOxZeKfLX
tFGx36G/e7438uOC9Z51xkbrQlMz6RA7HeLklle3QFfWNQ/XgMarIrA5+rqArqNr
KUAdo5/Mws7Ef5G8INk6RjMQdte05eVjr33qHfgS4q/Fy9rIbuDbZo4XvNWZnku6
n2pklAow4x3BRhurzSZPp/XWmWnRgu33RwWeZS+cAEnyk04aoQJ7YuH4DVazUyjJ
qFU/icBoJvJQXnvQZyfegB+14UgfM4koLOFAp9k+PTD//+gd1abf615sOIgKROdQ
LRvWvBhHUi5bZI3TwJuGtw2nYIWjbHNJaN2MlwP1W23fDe73a7uA8zWNbwZ0wVFH
RtrqVL8+DpAzMWuSMIpC1/5JvOlMLUjEw5A6GruS3rueDETEbt2RmfLqS6Ui3hcT
hMUrxG/Id5+UZrPrz/RFHZiIPG2st/G6a3/CaZCrbVH0nW4/Id/lI0yt1x88nSJq
95R8AUapqZuZyuRnKGKevf6L6rEGsmjTJttunchR7EsklV14pXVzk8Z5FwrDaD4V
r8G2kJiDn/G5s+ikqZ6VZs/8XtgWJKrGyROKuxF5sIcJKKFIFd1nprvQuJpLSkZc
SmLUsYRtbtmPsF9+/WUTstnWnVDfStzXlFMEHHgM6rTaialQsRLA2GmWiUYycaOm
0Xw4iM+pGv4ZTATYv8vfAsvriC4UxuIeQaLUHXm/Z7L19U7WfiB4NyGyqadMe26X
k5T/KzXpD1sTbFt3W08TJV5gJ3XAioXFPCvkhBy9jd6912gX1e1B+C5+KD6ZqZVW
K9rSxMLhCQyMmg79VUlILXZLToVrBY7TnqCfuJOFBt3D4anUJ8n3sDt4GeQVyWa4
9/awkbEkposI75KDf7tStoeNL8siLlw0dI/0gLPP+NFmGJadSfEMGpbnTUzXWUqs
sidrjVOiwu7aeHYNbzTulAXcTtD1Tu/5QZHcPdpADzaREVlXN7AuA9q87VpVwQsN
LK1T2yEN+pQqTiNTrksbdPlsPYZMUokkp5fGJdgG8C/UKEBZhujoWhYIRwY6ltEn
6f1IwInjdGKVvj+ULwph3ay8nE7pMrPCTszSNgUvTRF9wR3DCf1mE9fcGerXO8FN
LZXhVSILTHlo0gLtnSdV11DxoEt5yteisFzIlU5uDccVLwhb8QXzeIKe0+n3fwAj
cpFaRLrl2SW5KZJ642TloxVxgKNX/loQL1kJxmMusBoCDNE6hWoRXaLf1356oxSC
uaasrQdGyd+KNraRx35uZYUq5NWTFEsdm6V+j6ajXQDtjWhCzZHdh3cT5r16qtt8
YdxqNTjyOirFxYOsYwGnRZ5kslgBoB2Y1Shydb6sZvHyZw41A/uAkibPYseIV2/y
PdwtPnYXmMuWXQAr3UJUXSZ5NQl/s6MSHoc6ipQ/S2qhL1OhjXDRgwlkbRAaLmZ4
nBrJA/3C9p0M81b8GdjMWVNQzYFpvB2z5R02RFobGtl/yQw5HGBCWOl4dMwDB7T6
hU4AEmAqhe5cHkU/g6nCtC3nIv6maEV2u6GGnGl3lZPQj+pLHEKSyj8LOsGk0rzc
J8xMRv441x4WE3hPdL2aSdhj+J/S3Tpy3JMcTBM9Aizl786EK1ryvil/2gSwnW2M
hQfqa3j+wbKqxcoy2ZBf+FTLtJSiUcA4tpQSlVY1Ef4E1+CDnl7xB5A9fPuFwPg4
Mit3+zK3gi0+v2FvPiXvm2LVq0RUoOQ2PfYmpwzlu+V1Qd6pYZgY9UIi7Ic3C8t4
jGRxW0pf2qktDCfgbcnYmnCNxu/iNdwbUY+47syPnFakzOAJghGsyLbFGLIyPKgT
SyDWCCcKlNwN5pkOAoZole3maQ1lVQ4QNcZK94+um6Ez2efCRLDcDdA2da6B6VnB
TvgkSB7bYGMbVIGif+++aBeDpRyogeSn2u/lfxONQfT2D3VmXJBJpHS7hMVCTh8r
mF4FKSpCLuxH8l0L0k3wC1XN7SW3UITzgwHXdsrzUGy4z+lR3MzIVBdDnH0rrf/+
11CXxYwmYU6/Er0+FlNfE5mtDAodgV7tyEydbhoNZD9I9NgygAIgMlMl7unqiEzn
HsOyFd4ixF6nkSKDqaXmei8w6gHId8VZVOrORHsUevuHpC1MWqCVT1gZip+phOJ1
8ixzeqTTVO6KW6OpMiseB/8jL8cAjtN/IkqW+iyLoSZCvfgK+wO1fX3+C+LsiNc5
XeNZJMqNu4AFiMYkxFWnN1LQxkpwfq5R9RK7dOOsAEx+3QNXoEWbkbI6WJXgOILL
33RItYqdduYpPSVPFxGO2Et2L4CiSjZVLrEvhsHIRnKxb4Asvum/IviaT1oqkTfz
E1nzlzEpf9/tbXMTStZDY52d/yuenyMXgs8Ox8p3xJDCKeE97MyBZ8fnDPW9plhj
nw9X+XAupwQ5vjXAn0mXF+N9KqL5CmxxdGEPa1PYeMxiu6QLE6XqWu+UiWnrP055
KmoxhRmUJqJWX4nM/D9EiqJpTip3AyRQjZqSysrAw8eeTvfPilUqP+hqx19+emEV
Rh6VCrakD2obIDLEtBIX0IpmjRckynggWkNojGloOq38gTAjTF8v+4DT956wUv1j
BGDoy28HO++CSKofZ0j9P7aBKoVoShSb25MNqywsPRNsdgVkJdMEIDQR2ZWdlFM/
r8LuPG5vasgJJY/w3kL4kTsTGsu2C1uSt43iUTr247iq1vireQnX9jc/2L/Hrf2b
B3tgFsHwSSjqBuyh+aez6m3nx4Jj7hiOqlD9GMx1k+jrD9zzXIALmzonTRWc9SIG
YnEaKYH83Hcl4EMOfJcT+vbB5woqS93E6C8Qn0yiIvpHk+eYYZkz0xL+P/GK3qX8
hOyo1TpVidvHKFdMAcjtoZCA9ZjD096q3eV97D+mpi1MFzXqlOZSS6xOQrf0S1kE
9dMa4omKIFAluCivpKg9O02ngDUJYvAH0evo3dzNNzxH5OhJZIZDQCw0nAAh4+bY
DwE7g/ug3y4tyyNvdE1RXLQ5XTL84dEhkuHbZjdFeTRWn/AgLjJsRC9n0i42Asad
p+umtC53HgrL0aZ0g0cuZiK1d5ZPW46IAu2OcWCkfnL3DACOAybKAcE13i/IZJNh
iduaIgu8omvk5HEP3wzXupxmnvwfo5hQsxfhbKTlEFGNccRPux+JFhDR6iJZzF4Q
h9/229zDwU9Q3IZKTEzwNomwYI9DHogSshk7ktnYOEgB7pBZgCVDr4hfT+1O/SAL
yDrN3ZtBSRJVuPWlwvHW1p89OTMwm6dXk4mCAa3NAlM4DwMMOoCTIW6tus7kLpxH
8Aj1zwlj3CnpsCjfbaH01GQMO/4TioFVwTdHFUHdU+1I6ACAJkmnmofq0WJu0LcU
mEhFt61CXBgq7aTbwuC9V1s1Fx9pUnoqDnuupVmoNzDnOAWwJcl5PeqhGt+iJN6/
K44njgyzAtJHxTK8At/en6qriJ7BF7NFNNJpJBZ2eoGrrevn32sm9eGMQH9Am2QT
EyxEIRtETW1hgzYMiH9eD/qEC7bP74g+sw3FUjuRJhN/q1Vuds150CA6q6ugCHfP
uHm53VFzfDl+xiq+CyEarCSMZq9GsT0gdOD8wnHCGeAKJEFhqtM2wam3rJSURRcL
5R+ZAYukdLtTNfQISRu7VA6uawu+6e7axkGsZfreSCu4oK9FE6TjL7mO71JEqP82
fd6ChPLfOu1EElAFmelfmbU4Aqy4B6c3y768izVxxQ6zEcdeMz8RaOjPP3KbLNBD
8ooOkBdHtWfW7NT7fF9QW4azT6+eLmR1e9zfdrv0oOSaJITKcKOyZXKMgICt0nxu
69qaMctgwr7RYdqCeNYMyjo35JM3a1fjBNj1m257XyT7kDn2G+3/10oC7pu+ovNL
MsNADlkWBIxSH0ocTL4MZvMqQH5mbPffztkPqLMUx8IstjHp0QIAaK0Kbda9vKh+
oJugyP4UsnSltOI4dMa6yYIKfn9ZZflm7MXJF4JNbJPKsDwO/dfEQqYTaBe9YLOo
01iNzqCP6+wG9425KLDlhFRrOZCkby0zWtdAF7aVkM8dN31nnI/McsBgW9YPOMlJ
kfV8pl3vrQv9h0NBaDaMA2lmkcsqp9DN1zRbib4BN8dLEFb4vt6EOcTXoV0nD5FI
uk64y8q74j+qMWWzeqVW3OaK3u9AXBR/xH8nvmXWmFO+sOgbc1olvR9ro453SEMU
azidcZC4orMxkRwW9F5BbS8LeeJ+RWpjjziUcushC5b7A9Ima/kqZJuRrj5qbI09
SxwroyQSZdhVZ+PdDTHYXSWRyZnfVaEX/9g9L/b/b8XMI/2/tT+K2JRlHb25gayw
XYSdc3v3gpA0BzHcq1urjw1xzgT5wO3LZQRk1VSxvKwBL8QENpT6XmmaPsaPtMAM
OZ5zDsm7ki1urPy3K4Dv5F6hnDQB6FuIcUtMAACH0RIHIpB7hmslCPwxBagVOCGv
9gr2FMX8K6EoRh885woD6uyRsj6rn3aUXT8K3bxpL6CUZIHg8AAY4qaUVgEQQuQj
ERiLeYo9XOKEuYi2LdDz+x6eSqW3hZaOvnsDTbZtK3AiYSjRMkrpHufKIhUiInmB
b+VH+U7gn/ABTU62SbNkBBPCCq99XS2jw1bh/dymO0/HgAv3lgPrJc4V3fEYdEHu
X/kvo2Lxvzh38wE0NE3HyWZKj5YhEl1Yzp0tAE3mTk4Rbh69W5zX3lhMwa/qgDdn
LsDhSoq3W4ls7A/LXgixUZmNBcwIUhfGen4DlfqRi/giD7Y6vIV3SX5b4w4DXZNw
NIuPbpGO1JwWA2sZkb3MCleDJtUmQ1zyElRoqHY3tWFEZBEaDF5+3K1lnB2Nq/+Y
bgdY/R3P6peX6Z3IT6nWpGgxmgaJA3WqChg2wbZyp2nQBCLJakj42R7//I0oq108
1PQ20PA3kDF3+MKo11iNurqYTzBpqpUbDBF5Q8IKU/u9zTWfpjyazxmLnJDEXFjR
fgzllLtIiQ73v7bk7JAlwqTSWOCZrU2YIQr82SeL2c++WVjoDp8oWPYRtyz3arcA
uMQ97Ohyo3SdM1L8+605BJlZQgyqSy/25LRO5ZnwuzjKka2N1DY7Kh8cI0yrzJpg
64wWMLLr+hk5ySYogP5D/27u5l/Voc4BDx+CWcJcnxbRO8xpL0r5gneGILWpBZS8
6vH3/NMP9pV9wHhWeAse6RWgnws1ABdIakQ4V9ba5ztIl2Vd8E4Cdea6TKPZ03co
CqS4Weip1NCESv3sTSavBSa4IbOwppFd074mk13Afsdv+bzcJtz/TqiwVCiYnzug
XVl3OQgaeRjr1HJDr3k2mnOAzTv4b32kv509lR44PfRdvyo1Ne9dcP3kwjPRvGTy
D+gEuq8lwoit5ztUqkMOcl/hq/CXdtYsqFzYhGS5I0rZc8y5vrcqkfGuJffLqUyy
QGn0tJqa90yBrNoOBRiivt5VIR7kZjPCuW55q3CwSZ+oqPO5OasESIgcMNpv7mm1
CfPtvBAR+2OoHmOGk7wgLv22OThs2BknWCXqrka/OvxieWcWSXxC8oLxU4xqJdYa
DTVnjhNoyBnq9ZQsUf5mfmWZC6B0/wb1zQAufP7QHyVKYKgGPpg6nVy7gmKrc3R9
lWQnVQoS73rLUkb8K6wXLfTbsmJRJJAv073EOwDtYhvqGe0tsZTAu6rX574STjt3
EzOCwZ8lZirlN9zviZcANMMGz2MEl0zf3c+0cREGJ5KVUdxxkiVQ1U6vQqR4qIkT
nRoOyNciJPbBj5aaJc4jBk9oYX5n3/hNmngq6sl7R93l2/atc+/+syVCGyx8c5fw
BJkCtYLAl8nes6MkiSQTQMZQDWkt6tuGRuIEpGJElnZ2zUFmrgTBu0Cv2UeQPrvb
QypDHS37JLHe6AZOnPruafb000727007KwY1a9Cy/M1uYU2IOydDYA+hi5P2DIU1
gICvViwUgP9WWFs3xcgYFBlFSK/jXVzcWJ4MlHTOzNyD8tpaMhecrMEuB5VEqL3+
rMYeCrKR6Qvl1jvjvSOBroBXx9XOAx2qFU0vQ+iwn1eEb0kppaYg4gQEdTVDU+FM
QChbFMr30p2izjE8MDikrD51R4kXYdUfxG8q9XPP0tTPS4RPUs2zQRG1seAd/trH
tgzY+owFg6UnGTj85RYV8+bMNNG+CPqawFX1v37dzw3AbCAqp3JcObvdv5NRfvak
dFGqrGMIioJriX/UVMqIEIj1+9m76dfMHQDB9pdu3IsPQKkajPgqMA54wDn9VM/C
l6HHWKbII7aPsyxi1LTiUqk0ibOvka9Xc6Bj+C9EmGKDnXwKIhOXrMvb8w6wcmEu
QfvzWOF7q5JfBql1Y875wPTCZw2k3SlCB+hizsUpPxZ17U76ESXYe4aaoAvGVQfY
Af3rMuDehWA484uOjBRNqj+4WalacCJnwOjGwroKgybpZPbaS2SZB0IR+lJnnhyf
0uyUtn23bcdlbsHHpI9YQKcwZj4dqUidZT4Md1urLtZYU6Q0E4ovK8PZ7uvmjlXo
lkoNQkp8vuq7Bfc5l/YsF0gIO+HV44SU4MAWurG77eEav/Xi691Dp9eJ6IhrWwws
4pFh+eHXlhPbm6+Nq3PMyFYWuenEqn8P1WNr7z9jRfD5nkmKobGDPa0kii8zwxAt
7XOJXtXVSss91FNTaKqhFaumC8nLE/b5Ip3YnC5lZ+j8Y1tJS2EBmfZNQBdHp88S
kV2kfT4ifQZEUvNJLpkq0meIOnB8wWa91chS+K7snvtWKRWQznr2PzGUCxk0LmCT
Il2/gfQD8zrw/QW3YnK0BUCB6cIR+QM0pa/Gt1jfiDpvgeTcCzCZiFdVeqq9+R9k
R60aHiZoInfHBk8hXewJxfn1washCm6/SEcgUNFoE1u6r/OlceVWOzunGQ3wgB8e
KGKPU9KPlAu9Vqkpg5IzrwpoW6QqGMac+CMPQNwK0uYz3IF3v6mBJBKF6TnSD56a
f6AhK6OvKjOp/oeh8y3FttYPUh4vL0FfNrFFhTOFFlkk6XdMRRV4c6YvcDN890Aj
PY457hDDyUh46p4ZpVTD5Tw0vsRl1sny3QRfucATfVMZmpVbP6MVixcBfLNz+BKa
YTg8waTZdhY0NE7UMm+x4+HQl3+P9IZjy/VLc64jFOWY5o+1ek1M2yngs1AmBp+z
JtkbN6OvBc3kBk9eFKVTpkPncqD+E/dUoy0wyim0kZqJJpRQbL9j5hg5PXzf+hn3
DNhszUN9h02Wo2EZoP4opU64Qt3Xv1vKNKUjYSi23CE1/RUzDwGiQcD4E7aFZM9x
IymM2VGqfktmlao9eBNvTiswN/i/IN22OHEsGQH+Z/DHXjxQgaXMFVVgDrI68Rkp
IkbwVKSXOa/6lVfEtNz1ESpLVeZeb3D2ba337bac3F+R1tgIN4qBm+z/p6bTT5Yv
bJsajLklHM5itt2cs6FztZGg5dQa2lVeuDep72kP3wGCwREbgKMP8IdJQDn/oE+V
U8s7VJ7U7C4vZIpJR0BVybK2IusET2w9LTmIKZM+Zx7tH2TI0bQJ6kxePTDxWaNV
r1UfZOQQMXquqDgGPvaatlM4eHbk13tHYqcizM9JV/9poZ4FYohLuswLnwvzQ9qE
AdkbxLf+ORrAXyqxL90c69ke8B8k+SqvlxNLAkxN11rol5QtWNgq1wYTXQdYuPmt
z4fD52U0suAdNPG4JuKOBgUyX1jplYTLjUDcTW/moUF4wqhKjQ3SxoWpJ+QOxA49
FPcXx+5QeSBRTu8/YdOFU3WIOlCVqPgAQu78DdkCS/Nj08zuicJKSC3oWV8v8vpN
u+zS9KSZhaYw5oZIByU+sZQdaR+kmRY5mpvpAi5n0CVrK+j1DbqaYwXDSJyOPIsJ
2jKg264IEtW3YzpPg8sej4r7KXCsscG1xzHJimPMcazX/2lWMMU/f1bYA0/saAHQ
TsaoliQa1dX0kmg+pRvlrJ60/4Q0UIPyN3YtFSuFz+c+OlU5iGLQvVrruQVezZxF
LCn/Yv8bUALRB5evufZK1quqsJ89j5vykbfm0XNenYUqq0OltwFaKVUqXfoIIvEe
MneR/I7o1evEV32QN/BlrruZI7SDMouQ32nfxj4TD1cEIPgAsQSDBXxVpg0JX7Si
7zSE6yBIleV/pXplWYnyFO6cyJ0nagGbbARox4PVUtfLABV4MxHBLwzaYeB1WmRo
aK2XOcA1W/TPBOtWXY9VBmnVk8ih+66/LlJ3RRx4DqEBZfl1ob2kAInbuoMTvASr
BYNB3oXVSMNJkg+2/KZJvM7KbGxi0jpwsBZInVXTRXoAO9B9ETMQ2bRfczO6+dBk
d0ndBQStv1yGZYnDOrz3aEBOMitjwswPokdEdMNzKG5K15KEpbmglvzetaAGS0zU
pqPBPMIvlscoGbzC3eDqVwdnylWwrQCLmVIp+zoOz3axUdmL2x/yi54kPNMVCAJ8
8puvi51kDq+gkih9Bg18ZrUR35PtDv5yOFtib5kKkz2afNeFTrNHumaRsbCNfRdm
yRUURF6PK6pMJ2qsW2pQNT8eSJ1swFXCuKYZuVl/brZVDdSVjl8taBjpJnP/grod
/xlPKdvv7ANNhoCkpcYHT53fQIHeYAD0W1AtkObPnu1NjDytZuiR0Y06hhNKyn4J
5E4hhA5EVfHgVblYWeTmB+8AzV525Qw8rrZVIT3rQa4qoRJnk8JKPq1C4cD4cKD3
mSG+quwTN2dPm5q44ADDzQF5cxumMFgQzfanUy80xQFzVMgjsYYYuG7dRpPWBGFp
w5vS8DLcaW0f2a2dYhdWs5uXlupo5nblxfwZ8eg/5UeVvpKM7jXq3xRiTefIkMjO
0z8tbaOyG2fQLI3Q3Jvr3kpnl6TIPoyldk6j4tb2pqx5BrLvLk28nYvbT5YIFB+j
w3S4t2Ir0Uwp5gBahlLFUSVfW0D3smEdONXuUhRGUmfYagkxUL6kYw7lM2gejJkT
/KRgoqubebOgSn+ExemrG46gkCCbqRE8vVuMAg/KEKanEWiQN2+/hrEKfNgGI128
PqHfyxxdOBdKRxe0TDVn2mZfnom6n1kBvymD3AeM3rU1nX/S1ucyKFqx1vyMGYVh
06SRWpNiSErnIqIcef1zOID1f8zzc/LBF+ISKR9ARqB6NFTKxNfMRnZLs3C9v1hP
Obv9LBCM2jDj/es23HJ2Nui2ZImTooDJWlLbEb+b/T7UtKwruFbUKlFi/oj6y4Qs
YoDmrwunxsOfvrw3pylIt/p6y7GhCAw4990oK5AB0L9KCrnr8jksBvILupfma6zA
9yj/lQzP2c6gPRg+yI9khstEyyEBs9LfJHcLp44f1A1sB0zy59FVxeMlylLFN0cM
Rb7iCEtEGFkfU7EW0I4WBq3tdN+Z+hgv2KldhimBvI+gb4Gdoer3+1H17yHCEGhL
XEirQ5FFJszj5XT6iEtVgZpXNOXVoIKhAz8BS9us8FMLsun2H9MnaYAVW5s36VnC
LIQhNm+OlfKdM55H1zyMWeEE9X3ICSLGHT+j2klCCvCU45HCTkUOWUTdpATzXxS4
j62JeQvK217I9ZXgs5BPGT6VtglDp0zG8pCgk4Hc2yYaYNAICPQ2YfEVDWGMEDYv
LX75ffrWYRcBvpcgmfgtjcEsaoJYOY4PxX4E5tfz+S0fISwFcyMWH8nS3U2eNnJR
sbtZi6sDLTM3K4eNIUyBEqpDbZB3I6v5vTaHEHw+2otCsraxWhG4cxU828tUTmob
tAIjYMlC3i3HdtX9cXQ+mJRe7296jkLU7lzs39IuFzUshlottMb+bemT/Dq8a6Nv
PbC8ICbi2FrLku5w4p4pIXbmcONorldAmBpgqXgLh/7njzUk3l15DoN+4DpF/K9D
WSjQnXGItqCu0muY7If447kG6OB/l9//1LHURM3Huy3tU5A2PNlPrxeBIE2HcUbn
ggzfngZkUxrXNBKvIFRl8IxFwxtaCWl5XNBbh968FgLnhsNJYhmpQQddhbScAT5+
pn87j4YUXmJS8LUuS6sqsTS3TyRPG8Dv14Qq+g1OJn44inL9x5bL/9quZeKGQ+j+
JxJ4rj3aHB6Qz/VPl8ZcIFPFg3DV4p7kDAk0zSFAkApfsjnPkkHpyWclypoRrkQB
YJYCZvtX5WczUPxL96U3nLfjyPsFh8hgaVX/S673D4Qsk3wFXN1a6/iCYjJf1XWr
ufxzyKs5i3jv4TZcwDj4Wwg4KxI71rf1hXJOaJNiiCmbsITPqi43JRkZnjs3i/GK
D/L9CRyZgPf1BBEQht8KUWH9H6G7fk5AM5g0u6zPqT/NoMEmL2F0vwREIOdVbAe5
sFxky+thi0UmcETiUuWRTf4LyWdmyLxj8KoFW1/+FZ3t+2NScDQmQtyJ/llQ+dJh
yCDApIzkTeDXL+8QyRyx8lAWZjF1SIvMuzuOybzxGps0O0G4T6HfnJhuEHRHUBIU
oX/PM+XZLvthb0QzUzOToXfMf+OGffIa+mt6EyZLHhu3H+6/sOKnThl1bN32ckdc
7ylPMRhoq158zwBz7qaJ+ec0SYkn+8q3lDq8+X8xqtxiQJ3XBJRFTu8wUlYbwqc2
lreCxRjdMiGOby97PrFlcroP9GO/9x2Z/BsJJv41AiGO0rt2kMS4o3Gf2hwcewz4
UKPplvPt4QYXKdEiKOAlkj3GZS+52Hh5XHLCkfU8AaRUEg7nekiRnQNRLV95RhMd
DwjrTQ2hLsFEQ67rv+gK70mlIl94BaPx32ez9TrwB/e0DZSXcBNo8w4p9VrvUUee
o9GgznRNejEoRhICX1GlYqahEXI+VkIaUYBRUKKat91c7nI6pqW6Qc0pQFE82PRf
05ZsigAw5wP2Phua3LM5hknbrwLEGH/aoh6QpEn4PlTj0h31KDkCHH+FpBN9hy86
wE0xbdUkKEz3us4ZYzXTub19vxo8IzaA00ihPDcQPtzgHWAiHg2zg4ew2r37uAZW
JyOk+K6oaotmRzNnQNSR/3gyxA3yVGrxH829S8hPeA/M3+gqFUB9LXxpRrYfM/a+
jlw7WKXs5GD/M6F3areh06W2DKpSn34SUWcGEiE4iId1mWzcLv24hEqmt9JPVfeS
yL1VMwJ/0Cbch4FCtFm+2y1BuDzwkKMo8JvMIjSReuy7O2+6r9j/DZMMIPQeunUm
42T9m7rCxLbpZcajJo79w7DalyyppwATBvmNpa8dPeTREKH8nkcEAGYrBPfxHmny
FLDNbZpJT4tUsuyVObPdfrQtDfLMWDLiYKHGuZmQ7ysTAzO0WmxgFOa/rGQ4BSp4
VYwsrNJhDsTW+WSSTaLpXnddFIJ8vsnROY2Yauw5DUsONe7yT4nHmRE6xOc2FcA5
gc11HAcQDefQ0mQ2BEhX7JYJ0Wbkdm33OMNsO3NvBYykA1JW3bfif0Ww3Vmx//QW
d5MNnbOHfQ890mGCoOWuE3dJrEer+kd7iw3OSBKyC04ydwPMkkGCNO4z7u5odF8b
CSKiyuf9q5cTQ4vVyUthIO7keIwY3XMpWSy/PkS71XN8PC8C9iOboBmWD+U//CQw
+QaSCNEU5IyLdENt/7r1emcVPkDVTw1OeZzfgPDxMdFV4ZlBk6vd6YIzn5MFfLrg
dbHSqZaLeslST2U33/8TBnK4iaBUWS9fTiwYDqwVBCf8eymaJg/Qi4QMkNad7YpZ
PamHy/Qs+vg3hf4qvPMzGSN6B/TOuc9HtCbIsN+0ZZnMnndnXSQzOtn7bRF5cfW/
CBcYKtVmlXSl/d3QkfWNviaUyavBY2ExyMzHZtZOYtBtPBZBswJRZvbZP3/WIK59
PVRRFrrFue8ZvEZ31mUuOu6gnwQ/pJXIhMRJRSscR8XSr6wqolIyv8+C3aECUbiP
+vc3RqDp6ss02An1cdpn+ye0IxxqysTw2yhGctTzO/O5OwbJTYCueZSEMXaupn66
sEI3tHlALxZeWolTAuMESLajRjYhbwvSE5Mhpi6zSLZEYuxfrhrGCdjyOuzkcSQ7
oRfXCMB73pWPRInAXFElDPKOOm5u8cwWEvUNjN8sFVdu1qigDbReZAnFXCpbeUye
NKrvyDJTOhsd8By9o0K2NV7fs5w0wcpBIwOy4Ij/9x+skPvjKE4nKWd9iUHIVHzp
jJboTLcwPW3UbHshTT3y6V2BJ4RLOgb2tMnjA5gKCVbjftf50LoYXdLgMF+wikw9
PQgoEuRZ+5s2Z6AG7oBvl/kb+l8ifpXaVOiL1vr+VYLi99T8X6am7wwO/DuyD0Su
EusDiADSIaV+fRWlRbpMmQfta9mZUb5gcxDFVAUzkpppBaM1wNCQRV27EbzXmtCW
B6zNmcm1Ps124fUg/93PIydeTx+Shr8NJRp5qyrgf1vFebGkJkCz2hL+b4Ey+Rb1
sZGHcscIYLUu0Bf3JlPanvT012RuXT+fNFTwiu+xxJEjkbCUhWei7Me7AfvJm27Q
05wkGDPZ6wd7sVObVpaAjSDUpCQHxkkuw3zYnc9Xqolf9wsc6M26TucytvHlpQ6P
HzeohBGi/QfUNPN/fvoC1V7EniTxSzrqns4NYGis0WjtIKx1nQ2d4E1I952BxnCH
cnYFelhrD3r1QIT83BSFXIGE+AA6fnShm7iD1fpOi/PZNx+oM71jDG7QFD8m8sEh
NrYygE9zwrH5LWpvEr2GlUvTRuodoLCDmXefxewcMmFCPEbmPIrFmZrfizoweSOO
erOb35oMjk1G1c23QTVsdFgqyLU0Rx2cwkM4QpsmjDtxp+yfcJSLGG8dynT9tNH2
hWrlOhNNQjjwpq8S3k8QAXuzxToAAdTZovaM8f7WNU+lG1cOmAxAIPFcnQAsLCFy
Tq36hEdj1881RKM6ASuoaSpaOvjuhdhn8oL19mDBUxspfcjcPY7BKL7HoZQYijtx
JAY0cS88ZL3rxOtkOm62EFtg+lyz88lCXhanzs3cWLrzbnz/vbCY82tSL4jK/yjg
dyoMHJnE0ZgA0pWymjhBDHf/MwP9BE9NnEr48WX62I+wxpyVfICsBWSVxhWqeUAr
4ToSBQoJX7aCvXFDv8DuyNF3B5LC2rema3GQf9nB2UcLKdpJvMgqWVfRf1E+c9GF
XItJ3+1lhFx4z9o83RNNZiYqqDt5UutSOHGM6V6SyV1IQY6xnxi6sezRrRhY1XwQ
OGX6x/0A59BfiF5+AknpmmJlB+GbVLijWZS9CfMr7l4ap8+jhqpReiTx5Du9BGku
tswvAs9x4+psCmJVfvlIY/cuERyoY9nvv+adVogRD75UNGpB8JLbCvS1n+dtJs/N
Bfpu7P/DQdDyS1YbpCS2PGHeyETspjobdpbccIwSjvgaROt6l7KZHL17ikElZMV4
byUvPE0cawFCA9KnrOqcnPGTVZGGhi+u2dyFf04RSSR5sPTKpbNNPRBWu6BgexXY
ekJAWjZQ2SZrp/P9y6tPpE4DG7COgly1TXFY9XPA1k3Vifb+6eG9WZE5p5gl0x/X
mUxLiACRHl0xCJ6PGUsrb6yhP+UxpBpZ9HgONDgk2i1HFegu3G8HDO9/j3RW5HOk
Z1YRBFZV1MVRP+IMaLKOC0KqQuZzhm+GCb4SyJtpTdEHVil3BAGt0fGW4jQMsa/b
Cl6EJ8/omr0e/46s4+bqRCBrX34fut+xEmIMRLYUlxDO8TMaqFclDGLVhgdz5p7h
U+QpCWPW8Lpo83svPTNugvwFaHsVkDYpl9Wtgscf/RfLDPU6U6+yKj8jQ/Cn+Yef
ZQZKBMOV4JuRg1eYG3nBFY0XmMML8mpZ5+OqPR/+Hq7vYuQiJaQlGo696outpIe8
l3jQ2xYObTjefAa2fC2LkOYp7dXBkOf+T3hg+94akS+iCRgG4lDooIzlI7daptBA
aK21blgLh9JkutCXhmFirNE0Dkw+DEK6wxgCBXbzLwQNMjyzp8oH3BTu92CYVSN+
EFjL0Jn1yT7+gO5zWA7Ri6T/ElKx+trMG4rprWlOZ3mr8BqATJ4zxsw9t/eneF3t
BDPHlcuOVcIsOG04uL9UADSml2zbTXh+YQdf+qv1mHS2SszE7/p0GhbkvCbW6viB
tb3+k+YA6YeeuFpC8sFh+P76vIY07v0l7FTLKwfdvNDvY2+45/cw5f48gnOjd9E4
PcthyKvI4lpgyx0wkj8d9cAUanzyTcz7rhW329jBrPG+jYQ+CrBCsn2Ovc5ettzh
EKgTFZU+suXnQU2YYRY7ThyOdny+TSS/KS6DeNCorm+bMzDbywElER2sm3xEpVph
spG1ACDBncQ78HiQg9WGwWMuHUZAj4aZIpQaqfZ2Rctz4uN4bWTJtcBRHr4YuFRZ
n/fP5gmR8YdwTepsgpd/cwkctm2eU2V0vTWe0Whb/iXw6SJYmCDqHtXlDdh0rK3Y
pu1wboI2UNuEjtNMUO5N/OqT9xuNsOLbwqk0MtX6FEmvReFvdAX81QRDzdvZCsg0
PXTNinofZ5rOAeptKNfTpiDDX2UtW1jVhvF7Hg8HQX+mcsQLpo3CI33istG8yBy6
YJkRSKGf8pkgCkMIKf4ZsZ6ItZCkYmc0hb9B3E35bNkOYfmGPuOGUfy/0fPeWac9
qegCVG4cMMmTEnVtjCszYYUUqhIT5zEkmv4CQ41FXnOnDddB2vZeCYffYrkt/iPH
4xYDJQYnV5XiHdynMV8VCNjEkclCypmqqejIYfchyB8xkfD4tRo4GnYbLpKPBURz
B32OZR0mXymK9I4uf2EzZeT5UC3m2qA+zUuFrdBPdAutVxTONLGosPHf2PL+qfiY
tgZPVby74mXgqH4WIz3oy/XFr5dfY+Z8jGeCTMqr/DjdxwDoj6TsX0fQ1JPpBksF
QzG5VHAxJ+hcMifaaZUlh39ZkYReyUght4r52mXX41dzJwZ9pPLG8GyNpyQWVVhD
eR2tjgn2c16Qu5Cu4DaFr2faddlNNnSYGAYvrLlIYHeVXblm/5WMicGA5PQcsdH/
pf6US/Pr19vc8i5J9hKLxM2LU9OdxHRoecNM82S++NaMv3jOH6nGD/GxykwcsQ1F
jMhWxWraaPrUzHS0zzb/Y2oZ3xKL7XoVFbBhw3JZxEYY64CQmUfMQSkfMsqBE4Fi
vMTTfCv6bM0DMOaOfr8rHXfmbB2KF66yYlyeoZsoVg/5eb3A4DCvabTDPqWuxK8v
Im0Ah65hhXQfN5+7gwzcKVQjfNDlyAxa4Ld3Ratje92eBUzUS1F14kYV6Q9PsJDI
9uFTVHDtGolM5vBdCk2cS2EmwMlcVQiYMJ/dyKZqjkaiZRysHqkIRhc520eOmV4M
oGzRW8ni+CfQ87tPa2Tbj2A4ry7lmWt5Md7Z/OMLrJFK2VxRZ36ctoFYk8D+MlIh
9hlDC1hlcponxpKC2unjb5BebHMFUwfEmIfcZI2dwqRr0cRbeRCR8S0q4uZ+frbF
VyOeR5Japi1XS3FHU91srQ4igHRkhSYFVvgaq3JVVNrf2wWVMKq0dKnKkcse6FZe
h6LUkA3rmdCiKGEJ80k5lpkWNT2lUI+UNXVMIhXi5otfEiTjmQouVRu32BgUviNx
WPfYQwCzlwC15zZd/OhYwz/iz6ZA7+o4OZlwtuzkr8iSYvp0znTQmm533PMcLgnk
kj3asfA/Td79yEaOXZ2FsdxlaysrMjY5a6Rkw2rUe3MQLl3Upx2HaRwH2rX2cCKc
pJ/MK103cwhOAm49uV8yET+LBrRHOHbqFMhf1qQQyHKDZyGAUUBRcW6r10K10Pbb
f4ulAhIl/Ph2ZXeYcUSGfQXHrI9l/AVbfk/PhPqEPynG7JwET9RMeIxnYXxumewz
mLyZ+vPSXAQqhKB+V13416r/n1JQYYAPM8NxEhunL5JXmSrfnBZTDrfTRlCNBuDq
SK3YoX1BA57bPP0/K0HWr2sldtF4RZNLYuslwBD5jPV8RvHw0Auh0AtwGS/8UPTI
P65pqMvJoVk5WiJcI5Yat88ELd+aGhdki+6jq3+JqMX52c6GY3KdsoVCyqIFyPCo
Ks6esx4DDrsXk9r8jdhzArhqHWu/bYxveF0g9UHq5S0GKOxhXKZzrsMkI8SbBYRB
vIU1jCd5SW6ecKELs/VElyvv4X/Cvnju3S8yYwWnIEVl5O7oP+6GuvkejOENIiBR
TLVPVkClYBQmmGo4uI2K95/an5lLsbrotvcKHg1sbVkORZt9KSK2KmzYfhFF4t+y
qvVR4TB+1ir+4efMlRra/jq1IaKxEj4LjcayaGmfwx+U6rizp5HK5UiIEli7ZeRH
NXSLaskZaSiuTFs4r25jXnDV/aqmTcMA/eCc1d7B5U/oRQpHryngqtSM6NJg2Zlk
ng0RGk8Pl3At4aXKZ/fkf2MTLXa9cPp2Ae/Ye95NsUh80Gh4iVmQiFpGCvGYPrOh
OV8P9pg/79+0+4BHvrd9ifpqnrj2uOhfJV4MDrhe+HWdFCFwzMJ2Vc2SFItcd74r
mIufpi7JgzRYZIoI6/+k7J1vT8W3uwTuqB2DfEGubhtk4FKRJWWhinPbKdJpYhdU
CtKHGGfpMGd/Zg9jhVgmMpNXdU2vzEKujtEm9/MAB/0B3sTq0BeqCIhkIMRuq8CF
sKo/HVYgLo/Bo8bqqPd3vIkLsG06yBSBCMQO2jPMsNZ5vYDpQFUhoL7xl+xN3NPw
xUV3aUvKzcFSLJcNZK4ruwTdf7dBKrSYkkeBKCnKpi72qTMTY6aNiKeqYWdhwXfT
zrKUEGh1LTl8iiyMMc1ypVABXsMYFn/QDnbunahkjqh2BDkRpVnCmUBCPUx2ld4g
XxWU+82jzaCisSf1upvwDSZ1Bpyh94BUPvw7xOA0BcsUtQhSidW4zUneW4HmMwDN
ZJQwkqPYsYP5GLeOijJC8EDOXNNIDki2sqhNgcsKcyeGrVhuy1yjKYKPAG+C9k2x
I5v0MzAiOasyi5lBjdYFUg4ekTdj6mxliVTqePJvVBIcDcRHWX1tuOiFmk26Q4K+
BYugKXmpsxFTD+ZyinmdrMBL7zyjCmZSUWfzbv9AOTB8MVWR18vVJMfNcgUGOM0h
4rdBufU2QkHQSWqtWBjgjJT+zeRe9EWJ5DCLZJssRx6bRuhj6XU46ukxHJQrX9ie
mCq2b4IuoZitaoAfIsJA0aj0eT6k6zzd4s1EjL9ghSNMX7YXKgv6GT/Q+UPnQhWa
ERAihsxnWDYFrMkzCGe8SytRkR0AXsSeTwMcGXCJj/APZWPu8jr6ycZwcD2h5VKJ
ABM8MhrRbD6yHjOL9h1O1yh5qonFmMBfSsl+nfBe9rQdV9YG5ez2g1yZILnQH9qy
Vyb+nMc2GANWgAzQOLQMZfJkVcHkJVFdmP5bKr4Xnm579JBDSRmJTy4IaDfaDrAZ
fcXptLIDrWG4ttmK77KkHf/nOaODS6KeYgCi+GpHbjxVx4DO/aFOEJf1dDlm69yO
gQzhnk5kDnSWDDR6R3JEUz5dIL4Ex+dyU3cKC/2l8U5CcaQA61mSqeaPKczQPnaS
xEwwyaMdAABMXbme3CpRWcfAwi7wO2DuntdzvjvPN51DcNSAXmmH89lAeL9bQlCX
fSTiZZ/hfunYp5zHKou3gdg8Y7HXVPamokqkTraidxZlyVbacLp/7GSNBFTPtxJz
Pj43NI754pgc8I1t0fR5v3OJvKYJb8o6ANOpWEnsHxYX6ExK1uHuF46hGZ+4IrGU
B2MeSa9I8JH6mu7cc8prZ3uoTSXxN/abi8/1HGpTLevDmZqQHYfFjJSp2k0M3QX1
UkFYadsJti+u8toxScYUydrDCGb95a4v+bevebDYcP4a89n84ekW/YRWLe+bUisj
FgTioi0z2hdTUH5EXmqSuni8NB+NPsyelAaPoTBLILy+9cQeDLDWCPNszGbl4lQB
tLz3wFiGbYPtoyJRI9YuG9kRDASGqzW5DV+Re0EN2hGIA0Po7s97JPUumzPnUY0E
kQim4EB2m2KAl2iI/hEgBkix7AXRADPwLj6+YjL+0xG4BsApxKQxO39ziC8fJrhI
4AlBJkjOSx0+r+Nu9ksO2ekoAHVFd9ceaJNR0QKLykxyfye0pfkHM6uwEBm6unw5
VXhLFeRmiplXV+q8B7W1sJ87kZ/iZjwxCASymEdJGi/bPscVNDXJNhGbAiQ/igKr

//pragma protect end_data_block
//pragma protect digest_block
ni6q6ASxwDvODwFypNcTZq5k5G4=
//pragma protect end_digest_block
//pragma protect end_protected
