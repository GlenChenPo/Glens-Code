//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
eh3gDs31l2K9OPP3O/wum42RnvZntSaqvXnj/eD1xYlQkRhdx+wILMOM4k73WLve
W1iLLPA3nD9D0aIytyEc3WdMplrr1ShqS3eC/nVJ09z2wkT+PTtsMRUjPy9phA23
Epehz+TdP0b5ffuaTUODDscH6p3s4u/tWcCFR8PGsNA5t8KU47K2OQ==
//pragma protect end_key_block
//pragma protect digest_block
+7VsUiSHOmgYwBdzgkobvPvwNkE=
//pragma protect end_digest_block
//pragma protect data_block
91DNQo8h6E/sDcxTsbAyG8/IiUVkzG0762zHVNl0SJ2+sc6gag+hib5nQD0sc5pH
AG4s7mK0MUtusZFsr7IieJk03s4dIwqU83ngammrnAz7U9hv6r8hbthzxUlFAh/M
iJVW2T3+wCsotKxMlf0hsLJwKZPt2jwSPSigeyWQk1730sXr3M/IAvtUqpyr5bNJ
8d/11Je0pRvrqWgfrnJ9C/I33Xu30nXwfLT6XCoFjkA11HjMyqbe0gdk1OuDy4LU
2fJLVRnJmg8Af4Z07c0ANEqUepBaAhlCgqt1sgOEg8hAcCiHPjHspe+h13ZWQQG1
zUMgmDfDnLFzEhKZA+WvdQ==
//pragma protect end_data_block
//pragma protect digest_block
GY7KJVeY/lhUiUPYk4fIfaxtHhw=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ACbsfsqy6fA4sIJYzTPFboOv3N9StMwJ0wwWNBWVS/UANxiCbIrVZEhyMSITRYyb
8hFciDpzE6s4nlDspX06N9wY+frEG5Dgtu7FCxt36h89N+IVMSNIItVg0O9HY2lg
21RoHEa8098meuumdyPsd02Dk6+3WmKA2RPcjPd8hW+fIerKEF7eQg==
//pragma protect end_key_block
//pragma protect digest_block
mSn+Y0jKuAJRHH+OiBKRfZxXtdQ=
//pragma protect end_digest_block
//pragma protect data_block
wkEIGpm3mL2nb9eJ2dPp7hQwIQbvkHHd7TqHxxKQluydN0YGiwG9fULpFjXAlumP
96zLZIEdAk9qgfCdQApBaw0I8lc/nBzPkjB1scKa052sIuRzwCxS5AOCviZRnO3U
352xVDQxM3sUrLjximqNvSQnPCECZomKngAGNrF/7625hK48Vtz+xiqKwYq3Izje
h9CfvxLHLjKDEiq1A8IKBup2LgRsNJWImTzTav05edujEjgmgu2B0t5W7vaf+Gyg
HP7/OVIqdyof5VFvGtOOD6TY3WuhNRkiINsS6gFbnrjA9Oyg0mfaO97KSdV8oAUl
DRyDA7/UyAvgcItOg8S4ORZLn4NWVc9yilRCx6FsJYYUNhsPs/hWO0adX/6HXQPH
wAbZkmMdoStEyVhfHOyWRQeX0sV0d3eiNotZ/7pr7JEL+vXXKhIED2Y8pptN0OYE
Qvy7zbn1YOQB2OEYnd/SZU/Pi+nNfof9WH2y8O5AvtrfyirOo76GyBhfRfeiZcMP
jbePlju0zpltMOzVGYCtGdFZqmm6kjMgmg6RoojoSgr2YPmW+eqRnhYru+3p2X4q
9sHhQvrns/s+yj4FsJ9YJ5CWI/RSom3hV0ncO7fx2sEdSJ4I1wRH+PvprTp65vQr
oX5489aKRaWxIAvfF/L71K4yWCnRQLpqq9Oevmj/Mvj32jSWYkyl7Hd1bkH4Yd8+
8H2e4lOLIWvExRD4qMDzmVp5jG74cVTICku6DK8cb2gZ2hxu3mWkQuCgbqfVhs3u
CEpFdWWpCrOe4up3BmVXTNktmKKgF0ztwMsgSR2X2jc1BHO/sji/aT4kjfLIM0qa
3XmC7l2iWunLYDHixsPJ4QRZUUL1ZZ3WhlzZQhYH/6kMW3UOwn93A/E6jlJcP2fY
xfTlx2STnYT+QAg3i47KhABvL1oSiLDw6UkiCuiBg1eYxUZbag98paE4gaFP7KzF
NgYL/LIWmEvRaBKbOWJX8KPer44bnvok32mFctHEWEKUE2witoy3TSgOsM+qAX+a
NLUMqFSLfib37aiGCRNK/WRtWEKMXXudFa48GDFttHVa4D1weTEpYcQz/Oj4Thoi
N2cNAv2uE4T7qRz9vbnz51lX7UH1gW8cQH0fFR62NzxlKhBNwCJIjOaE/GgmtER6
cBBIw7s5PxYlvzqCX9ocZJ9BZ2eZs/a2qmfQhk+yk8Y76lUe7VulppD1P8/zhlYu
xrgL8iNPpVdENTg6thyixTkkbPb6wbTM9eFto7RqJW+lUCP7V9xCtkVXt8+5r1eA
kYo7hZ8hssSEdGfLFQMMMItQrf/uIHoXE7HVkT4BcMYD4Bkz82bZ4jdRjaS67gLM
3isBU40+WrztDQWcHWuJCmbUarg8Ez86fu8s8fty67V6FYDcEuJeDdVYVN6bkiuz
aDj92j3v27lmuoowED9q3zeBWKY+gzY9lb3mLB597qov1JvuDFLKOkom22MnaTJW
iXotS4rVNLuK4BYr3QtzeFZHt1MoNpfZoo7kXHcIAHjrUoeFVJki9/Kd8uOsdJZk
Y4cxkItktb1z8uk+yVdBjfwPUezaVwFhNDOu2GGVwAdeQkMYOjsumvG3CClRrcas
H6rpRiy5zuXih2ZAWPqZpKyBRQ1NPjHf4tSOwheQiLKk7cfkbbiYRifBjalsTSrD
Ez2BZ0CWL713kzUfGAnJNVOFdMcJeQBNEu3I+iJ5f3ODX4AkUtc/yVLtuxuo/PWi
ilS1477tCRxVw3kkTaFydVVv7r2pRaSjXNyuXM36PG4zuQ3k2KL15247gofRSEFg
Qf3m407REvfvejXo7Icl4o4BVlkmFNnzSrIMUX9vVl6yQxJkXaQoW0pXqRA1zLaz
88ThG1PTJCwxdem7KaUtrBHy1JDN5PmONxIIPfCnOJJSsR9cuTJc33j0X8vPeh4q
VjizGAzCCKuvILVDDESvxHwuJof2+kVMlFg5ZzL64NCN83MPWh4HvDQ98/AbPIgP
jQBTgy5F2lAaK6NdG88pVVHRRGjIq/2GdntWJM46FFyIjGUG4krnsvnGkdHmJjjl
gU0qXB4u+TMrfJUyNlpp7cM3TX7XDTA+rmmK9V2oMZ5P5Iw4KgxvzWNYQuC1a3+D
KHKyySZOwNPyL9Ob+KxRdMqyCs/ykAqPM7PfOC00O57H0zXnlkhf/1dFr+7t/8e1
wEKm4n4eX+ihaWs81yH5GvAFqMRmVOVrVkP+sLO4FLyvnPKLiryKw5WBeBPI23yi
mb87VHg4RSHsoXu5zi19I4Kf4LX59BJodoTJt5UjS1hDZMwot3zPxZlYbTSuwm+h
7PaWHGNim14HvUGImE/NSzSFgATQ1rTCGv3NuZ/MigWxxZ8mdTA/N/mUW8AeE9mn
7cwHrYWKQ9M6Pza7Zu7kqoVVAd3e1lrplCJvamWbCtTxiNxSJZidXN0IYSld27Oc
w+OD/QWGTeMfHtVOEQI97eWueQU38w6NLedFL11UlX8j2Nxrlmz8mml/zX+/Bcdn
2dhHLwnPotAivZLcep6e27UP4rP5d33FMLdKs3MJfUrJ0lxtQ5atqrf29Scwt7+i
aj9mpGIpYNiamdHPZaHVbw==
//pragma protect end_data_block
//pragma protect digest_block
Dlt6kvOioR7pQrUvbGPNkQ23lOA=
//pragma protect end_digest_block
//pragma protect end_protected
