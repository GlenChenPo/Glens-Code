//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   File Name   : WD.v
//   Module Name : WD
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module WD(
    // Input signals
    clk,
    rst_n,
    in_valid,
    keyboard,
    answer,
    weight,
    match_target,
    // Output signals
    out_valid,
    result,
    out_value
  );
  // ===============================================================
  // Input & Output Declaration
  // ===============================================================
  input clk, rst_n, in_valid;
  input [4:0] keyboard, answer;
  input [3:0] weight;
  input [2:0] match_target;
  output reg out_valid;
  output reg [4:0]  result;
  output reg [10:0] out_value;
  // ===============================================================
  // ===============================================================
  // ===============================================================
  // Genvar & Parameters & Integer Declaration
  // ===============================================================
  // state
  parameter IDLE    = 2'd0;
  parameter STATE_1 = 2'd1; //get the input
  parameter STATE_2 = 2'd2; //process
  parameter STATE_3 = 2'd3; //output
  //genvar

  // ===============================================================
  // Wire & Reg Declaration
  // ===============================================================

  reg [1:0] current_state,next_state;//current & next state
  reg  a0,a1,a2,a3,a4;
  reg  b0,b1,b2,b3,b4;
  reg [2:0] A,B;
  reg [12:0] cnt;//counter

  // temporary
  reg [4:0] key_tmp [0:7];
  reg [4:0] ans_tmp [0:4];
  reg [3:0] wei_tmp [0:4];
  reg [2:0] tar_tmp [0:1];

  //reg [4:0] sp_wei [0:4];

  reg [10:0] val_tmp;
  reg [4:0] cmp [0:4];
  reg [4:0] cmp1 [0:4];
  reg [4:0] cmp2 [0:4];
  reg [4:0] cmp3 [0:4];
  reg [4:0] cmp4 [0:4];

  // ===============================================================
  // Finite State Machine
  // ===============================================================
  /*      cccccccccc                             cccccccccc
        ccc   c    ccc                         ccc   c    ccc                                  
       cc     c      cc                       cc     c      cc                               
      ccc     c      ccc                     ccc     c      ccc                             
       cc      c     cc                       cc      c     cc                               
        ccc      c ccc                         ccc      c ccc                  
          cccccccccc                             cccccccccc                                       
  */
  // -----------------Set Counter-----------------------------------
  always @(posedge clk or negedge rst_n) //cnt
  begin
    //Reset--------------------------------------
    if(~rst_n)
    begin
      cnt <= 0;
    end
    else if(in_valid && cnt==7)
    begin
      cnt <= 0;
    end
    else if (cnt==6727)
    begin
      cnt <= 0;
    end
    else if (current_state==IDLE && cnt==5)//cnt = output cycle
    begin
      cnt  <= 0;
    end
    //count-------------------------------------
    else if(in_valid)
    begin
      cnt <= cnt+1;
    end
    else if (current_state == STATE_2)
    begin
      cnt <= cnt+1;
    end
    else if (current_state == STATE_3)
    begin
      cnt <= cnt+1;
    end
    else if (out_valid)
    begin
      cnt <= cnt+1;
    end
  end


  // ----------------------Current State----------------------------
  //----------------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if (!rst_n) // rst_n=0(idle)  rst_n=1(next state)
      current_state <= IDLE;
    else
      current_state <= next_state;
  end
  //---------------------- Next State-------------------------------
  //----------------------------------------------------------------
  always @(*)
  begin
    case (current_state) //Current_state
      IDLE:
      begin
        if (in_valid)
          next_state = STATE_1;
        else
          next_state = IDLE;
      end
      STATE_1: //GET THE INPUT
      begin
        if (~in_valid)
          next_state = STATE_2;
        else
          next_state = STATE_1;
      end

      STATE_2: //PROCESS
        if (cnt==6727)
          next_state = STATE_3;
        else
          next_state = STATE_2;

      STATE_3: //GET THE OUPUT
        if(cnt==4)
          next_state = IDLE;
        else
          next_state = STATE_3;

      default:
        next_state = IDLE;
    endcase
  end
  //----------------------- Output Logic----------------------------
  //----------------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if (!rst_n)
      out_valid <= 0;
    else if (current_state == STATE_3)
      out_valid <= 1;
    else if (current_state==STATE_1)
      out_valid <= 0;
    else if (current_state==STATE_2)
      out_valid <= 0;
    else if (current_state==IDLE)
      out_valid <= 0;

  end
  // ===============================================================
  /*    SSSSSS     TTTTTTTTTT      AA           11
      SS               TT         A  A         111                                              
      SS               TT        AA  AA       1111                                                  
        SSSSSS         TT       AAAAAAAA        11                          
              SS       TT       AA    AA        11                                                 
              SS       TT      AA      AA       11                          
       SSSSSSS         TT      AA      AA    1111111                            
  */
  // ===============================================================
  // proc_1 Store the keyboard
  //-------------------------------------------------

  always @(posedge clk or negedge rst_n)
  begin : proc_1
    if(~rst_n)
    begin
      key_tmp[0] <= 0;
      key_tmp[1] <= 0;
      key_tmp[2] <= 0;
      key_tmp[3] <= 0;
      key_tmp[4] <= 0;
      key_tmp[5] <= 0;
      key_tmp[6] <= 0;
    end
    else if(in_valid && cnt<8)
    begin
      key_tmp[0] <= key_tmp[1];
      key_tmp[1] <= key_tmp[2];
      key_tmp[2] <= key_tmp[3];
      key_tmp[3] <= key_tmp[4];
      key_tmp[4] <= key_tmp[5];
      key_tmp[5] <= key_tmp[6];
      key_tmp[6] <= key_tmp[7];
      key_tmp[7] <= keyboard;
    end
  end
  //-------------------------------------------------
  // proc_2 Store the anwser & weight
  //-------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin : proc_2
    if(~rst_n)
    begin
      ans_tmp[0] <= 0;
      ans_tmp[1] <= 0;
      ans_tmp[2] <= 0;
      ans_tmp[3] <= 0;
      ans_tmp[4] <= 0;
    end
    else if(in_valid && cnt<5)
    begin
      ans_tmp[0] <= ans_tmp[1];
      ans_tmp[1] <= ans_tmp[2];
      ans_tmp[2] <= ans_tmp[3];
      ans_tmp[3] <= ans_tmp[4];
      ans_tmp[4] <= answer;
    end
  end
  //-------------------------------------------------
  // proc_3 Store the weight
  //-------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin : proc_3
    if(~rst_n)
    begin
      wei_tmp[0] <= 0;
      wei_tmp[1] <= 0;
      wei_tmp[2] <= 0;
      wei_tmp[3] <= 0;
      wei_tmp[4] <= 0;
    end
    else if(in_valid && cnt<5)
    begin
      wei_tmp[0] <= wei_tmp[1];
      wei_tmp[1] <= wei_tmp[2];
      wei_tmp[2] <= wei_tmp[3];
      wei_tmp[3] <= wei_tmp[4];
      wei_tmp[4] <= weight;
    end
  end

  //-------------------------------------------------
  // proc_4 Store the match_target (_A,_B)
  //-------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin : proc_4
    if(~rst_n)
    begin
      tar_tmp[0] <= 0;
      tar_tmp[1] <= 0;
    end
    else if(in_valid && cnt<2)
    begin
      tar_tmp[0] <= tar_tmp[1];
      tar_tmp[1] <= match_target;
    end
  end
  // ===============================================================
  /*    SSSSSS     TTTTTTTTTT      AA          222222222
      SS               TT         A  A        22       22                                           
      SS               TT        AA  AA                22                                            
        SSSSSS         TT       AAAAAAAA              22                      
              SS       TT       AA    AA           222                                                 
              SS       TT      AA      AA        222                            
       SSSSSSS         TT      AA      AA     222222222222                              
  */
  // ===============================================================
  // determine how many A&B cmp[0 1 2 3 4] have.
  // ---------------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      a0<= 0;
      b0<= 0;
    end
    else
    begin
      if (cmp[0]==ans_tmp[0])
      begin
        a0<=1;
        b0<=0;
      end
      else if (cmp[0]==ans_tmp[1]||cmp[0]==ans_tmp[2]||cmp[0]==ans_tmp[3]||cmp[0]==ans_tmp[4])
      begin
        b0<=1;
        a0<=0;
      end
      else
      begin
        a0<=0;
        b0<=0;
      end
    end
  end
  //---------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      a1 <= 0;
      b1 <= 0;
    end
    else
    begin
      if (cmp[1]==ans_tmp[1])
      begin
        a1<=1;
        b1<=0;
      end
      else if (cmp[1]==ans_tmp[0]||cmp[1]==ans_tmp[2]||cmp[1]==ans_tmp[3]||cmp[1]==ans_tmp[4])
      begin
        b1<=1;
        a1<=0;
      end
      else
      begin
        a1<=0;
        b1<=0;
      end
    end
  end//--------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      a2 <= 0;
      b2 <= 0;
    end
    else
    begin
      if (cmp[2]==ans_tmp[2])
      begin
        a2<=1;
        b2<=0;
      end
      else if (cmp[2]==ans_tmp[0]||cmp[2]==ans_tmp[1]||cmp[2]==ans_tmp[3]||cmp[2]==ans_tmp[4])
      begin
        b2<=1;
        a2<=0;
      end
      else
      begin
        a2<=0;
        b2<=0;
      end
    end
  end//-------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      a3 <= 0;
      b3 <= 0;
    end
    else
    begin
      if (cmp[3]==ans_tmp[3])
      begin
        a3<=1;
        b3<=0;
      end
      else if (cmp[3]==ans_tmp[0]||cmp[3]==ans_tmp[1]||cmp[3]==ans_tmp[2]||cmp[3]==ans_tmp[4])
      begin
        b3<=1;
        a3<=0;
      end
      else
      begin
        a3<=0;
        b3<=0;
      end
    end
  end//--------------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      a4 <= 0;
      b4 <= 0;
    end
    else
    begin
      if (cmp[4]==ans_tmp[4])
      begin
        a4<=1;
        b4<=0;
      end
      else if (cmp[4]==ans_tmp[0]||cmp[4]==ans_tmp[1]||cmp[4]==ans_tmp[2]||cmp[4]==ans_tmp[3])
      begin
        b4<=1;
        a4<=0;
      end
      else
      begin
        a4<=0;
        b4<=0;
      end
    end
  end
  // ===============================================================
  // compare the AB==AB
  // ---------------------------------------------------------------
  always @(posedge clk or negedge rst_n)
    if(~rst_n)
    begin
      cmp2[0]<=0;
      cmp2[1]<=0;
      cmp2[2]<=0;
      cmp2[3]<=0;
      cmp2[4]<=0;
      A<=0;
      B<=0;
    end
    else
    begin
      if (current_state==STATE_1)
      begin
        cmp2[0]<=0;
        cmp2[1]<=0;
        cmp2[2]<=0;
        cmp2[3]<=0;
        cmp2[4]<=0;
        A<=0;
        B<=0;
      end
      else
        if (current_state==STATE_2)
        begin
          A<=a0+a1+a2+a3+a4;
          B<=b0+b1+b2+b3+b4;
          cmp2[0]<=cmp1[0];
          cmp2[1]<=cmp1[1];
          cmp2[2]<=cmp1[2];
          cmp2[3]<=cmp1[3];
          cmp2[4]<=cmp1[4];
        end
    end

  always @(posedge clk or negedge rst_n)
  begin
    if (~rst_n)
    begin
      cmp3[0]<=0;
      cmp3[1]<=0;
      cmp3[2]<=0;
      cmp3[3]<=0;
      cmp3[4]<=0;
    end
    else
    begin
      if (current_state==STATE_1)
      begin
        cmp3[0]<=0;
        cmp3[1]<=0;
        cmp3[2]<=0;
        cmp3[3]<=0;
        cmp3[4]<=0;
      end
      else if((A==tar_tmp[0]) && (B==tar_tmp[1]))
      begin
        cmp3[0]<=cmp2[0];
        cmp3[1]<=cmp2[1];
        cmp3[2]<=cmp2[2];
        cmp3[3]<=cmp2[3];
        cmp3[4]<=cmp2[4];
      end
      else
      begin
        cmp3[0]<=cmp3[0];
        cmp3[1]<=cmp3[1];
        cmp3[2]<=cmp3[2];
        cmp3[3]<=cmp3[3];
        cmp3[4]<=cmp3[4];
      end
    end
  end



  /* =========================================================================================
         if it is bigger one that we store it to cmp4.           *****************************
                                                        ************************************** 
                                                  ********************************************
   ------------------------------------------*************************************************
  */
  always @(posedge clk or negedge rst_n)
  begin
    if (~rst_n)
    begin
      cmp4[0]<=0;
      cmp4[1]<=0;
      cmp4[2]<=0;
      cmp4[3]<=0;
      cmp4[4]<=0;
      val_tmp<=0;
    end
    else
    begin
      if (current_state==STATE_1)
      begin
        cmp4[0]<=0;
        cmp4[1]<=0;
        cmp4[2]<=0;
        cmp4[3]<=0;
        cmp4[4]<=0;
        val_tmp<=0;
      end
      else if (current_state==STATE_2)
      begin

        if (cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4]
            >val_tmp)
        begin
          val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
          cmp4[0]<=cmp3[0];
          cmp4[1]<=cmp3[1];
          cmp4[2]<=cmp3[2];
          cmp4[3]<=cmp3[3];
          cmp4[4]<=cmp3[4];
        end
        else if (cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4]
                 ==val_tmp)
        begin
          if (cmp3[0]*16+cmp3[1]*8+cmp3[2]*4+cmp3[3]*2+cmp3[4]>
              cmp4[0]*16+cmp4[1]*8+cmp4[2]*4+cmp4[3]*2+cmp4[4])
          begin
            val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
            cmp4[0]<=cmp3[0];
            cmp4[1]<=cmp3[1];
            cmp4[2]<=cmp3[2];
            cmp4[3]<=cmp3[3];
            cmp4[4]<=cmp3[4];
          end
          else if (cmp3[0]*16+cmp3[1]*8+cmp3[2]*4+cmp3[3]*2+cmp3[4]==
                   cmp4[0]*16+cmp4[1]*8+cmp4[2]*4+cmp4[3]*2+cmp4[4])
          begin
            if (cmp3[0]<cmp4[0])
            begin
              val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
              cmp4[0]<=cmp3[0];
              cmp4[1]<=cmp3[1];
              cmp4[2]<=cmp3[2];
              cmp4[3]<=cmp3[3];
              cmp4[4]<=cmp3[4];
            end
            else if (cmp3[0]==cmp4[0])
            begin
              if (cmp3[1]<cmp4[1])
              begin
                val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
                cmp4[0]<=cmp3[0];
                cmp4[1]<=cmp3[1];
                cmp4[2]<=cmp3[2];
                cmp4[3]<=cmp3[3];
                cmp4[4]<=cmp3[4];
              end
              else if (cmp3[1]==cmp4[1])
              begin
                if (cmp3[2]<cmp4[2])
                begin
                  val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
                  cmp4[0]<=cmp3[0];
                  cmp4[1]<=cmp3[1];
                  cmp4[2]<=cmp3[2];
                  cmp4[3]<=cmp3[3];
                  cmp4[4]<=cmp3[4];
                end
                else if (cmp3[2]==cmp4[2])
                begin
                  if (cmp3[3]<cmp4[3])
                  begin
                    val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
                    cmp4[0]<=cmp3[0];
                    cmp4[1]<=cmp3[1];
                    cmp4[2]<=cmp3[2];
                    cmp4[3]<=cmp3[3];
                    cmp4[4]<=cmp3[4];
                  end
                  else if (cmp3[3]==cmp4[3])
                  begin
                    if (cmp3[4]<cmp4[4])
                    begin
                      val_tmp<=cmp3[0]*wei_tmp[0]+cmp3[1]*wei_tmp[1]+cmp3[2]*wei_tmp[2]+cmp3[3]*wei_tmp[3]+cmp3[4]*wei_tmp[4];
                      cmp4[0]<=cmp3[0];
                      cmp4[1]<=cmp3[1];
                      cmp4[2]<=cmp3[2];
                      cmp4[3]<=cmp3[3];
                      cmp4[4]<=cmp3[4];
                    end

                    else
                    begin
                      cmp4[0]<=cmp4[0];
                      cmp4[1]<=cmp4[1];
                      cmp4[2]<=cmp4[2];
                      cmp4[3]<=cmp4[3];
                      cmp4[4]<=cmp4[4];
                      val_tmp<=val_tmp;
                    end
                  end
                  else
                  begin
                    cmp4[0]<=cmp4[0];
                    cmp4[1]<=cmp4[1];
                    cmp4[2]<=cmp4[2];
                    cmp4[3]<=cmp4[3];
                    cmp4[4]<=cmp4[4];
                    val_tmp<=val_tmp;
                  end
                end
                else
                begin
                  cmp4[0]<=cmp4[0];
                  cmp4[1]<=cmp4[1];
                  cmp4[2]<=cmp4[2];
                  cmp4[3]<=cmp4[3];
                  cmp4[4]<=cmp4[4];
                  val_tmp<=val_tmp;
                end
              end
              else
              begin
                cmp4[0]<=cmp4[0];
                cmp4[1]<=cmp4[1];
                cmp4[2]<=cmp4[2];
                cmp4[3]<=cmp4[3];
                cmp4[4]<=cmp4[4];
                val_tmp<=val_tmp;
              end
            end
            else
            begin
              cmp4[0]<=cmp4[0];
              cmp4[1]<=cmp4[1];
              cmp4[2]<=cmp4[2];
              cmp4[3]<=cmp4[3];
              cmp4[4]<=cmp4[4];
              val_tmp<=val_tmp;
            end
          end
          else
          begin
            cmp4[0]<=cmp4[0];
            cmp4[1]<=cmp4[1];
            cmp4[2]<=cmp4[2];
            cmp4[3]<=cmp4[3];
            cmp4[4]<=cmp4[4];
            val_tmp<=val_tmp;
          end
        end
        else
        begin
          cmp4[0]<=cmp4[0];
          cmp4[1]<=cmp4[1];
          cmp4[2]<=cmp4[2];
          cmp4[3]<=cmp4[3];
          cmp4[4]<=cmp4[4];
          val_tmp<=val_tmp;
        end
      end
    end

  end
  // =======================================================
  /*    SSSSSS     TTTTTTTTTT      AA        33333333
      SS               TT         A  A      33      333                                       
      SS               TT        AA  AA              33                                        
        SSSSSS         TT       AAAAAAAA      3333333                 
              SS       TT       AA    AA            33                                         
              SS       TT      AA      AA   33      333                 
       SSSSSSS         TT      AA      AA    333333333                   
  */
  // =======================================================
  // Store score
  //-------------------------------------------------
  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      out_value<=0;
      result <=0;
    end
    else
    begin
      if (current_state == IDLE)
      begin
        out_value<=0;
        result <=0;
      end
      else if (current_state==STATE_1)
      begin
        out_value<=0;
        result <=0;
      end
      else if (current_state==STATE_3 && cnt<5)
      begin
        out_value <= val_tmp;
        result <= cmp4[cnt];
      end
    end
  end


  /*=================================================================================
          ccccc  cc cc  cc   pppppp                  ccccc  cc cc  cc   pppppp                                                   
        ccc      ccc  cc  c  pp   pp               ccc      ccc  cc  c  pp   pp                                            
        ccc      cc   c   c  pppppp                ccc      cc   c   c  pppppp                                             
         cccccc  cc   c   c  pp                     cccccc  cc   c   c  pp                                                  
  */
  always @(posedge clk or negedge rst_n)
  begin
    if (~rst_n)
    begin
      cmp1[0]<=0;
      cmp1[1]<=0;
      cmp1[2]<=0;
      cmp1[3]<=0;
      cmp1[4]<=0;
    end
    else
    begin
      if (current_state==STATE_1)
      begin
        cmp1[0]<=0;
        cmp1[1]<=0;
        cmp1[2]<=0;
        cmp1[3]<=0;
        cmp1[4]<=0;
      end
      else if (current_state==STATE_2)
      begin
        cmp1[0]<=cmp[0];
        cmp1[1]<=cmp[1];
        cmp1[2]<=cmp[2];
        cmp1[3]<=cmp[3];
        cmp1[4]<=cmp[4];
      end
    end
  end

  always @(posedge clk or negedge rst_n)
  begin
    if(~rst_n)
    begin
      cmp[0] <= 0;
      cmp[1] <= 0;
      cmp[2] <= 0;
      cmp[3] <= 0;
      cmp[4] <= 0;
    end
    else
      if (current_state==STATE_1)
      begin
        cmp[0] <= 0;
        cmp[1] <= 0;
        cmp[2] <= 0;
        cmp[3] <= 0;
        cmp[4] <= 0;
      end
      else if (current_state==STATE_2)
      begin
        case(cnt)
          0:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          7:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          8:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          9:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          10:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          11:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          12:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          13:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          14:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          15:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          16:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          17:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          18:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          19:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          20:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          21:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          22:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          23:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          24:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          25:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          26:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          27:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          28:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          29:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          30:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          31:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          32:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          33:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          34:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          35:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          36:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          37:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          38:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          39:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          40:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          41:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          42:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          43:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          44:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          45:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          46:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          47:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          48:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          49:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          50:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          51:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          52:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          53:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          54:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          55:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          56:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          57:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          58:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          59:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          60:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          61:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          62:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          63:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          64:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          65:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          66:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          67:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          68:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          69:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          70:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          71:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          72:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          73:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          74:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          75:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          76:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          77:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          78:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          79:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          80:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          81:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          82:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          83:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          84:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          85:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          86:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          87:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          88:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          89:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          90:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          91:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          92:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          93:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          94:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          95:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          96:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          97:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          98:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          99:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          100:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          101:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          102:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          103:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          104:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          105:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          106:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          107:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          108:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          109:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          110:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          111:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          112:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          113:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          114:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          115:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          116:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          117:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          118:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          119:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          120:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          121:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          122:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          123:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          124:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          125:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          126:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          127:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          128:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          129:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          130:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          131:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          132:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          133:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          134:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          135:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          136:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          137:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          138:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          139:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          140:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          141:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          142:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          143:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          144:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          145:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          146:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          147:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          148:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          149:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          150:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          151:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          152:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          153:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          154:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          155:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          156:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          157:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          158:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          159:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          160:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          161:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          162:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          163:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          164:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          165:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          166:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          167:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          168:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          169:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          170:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          171:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          172:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          173:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          174:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          175:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          176:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          177:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          178:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          179:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          180:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          181:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          182:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          183:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          184:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          185:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          186:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          187:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          188:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          189:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          190:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          191:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          192:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          193:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          194:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          195:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          196:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          197:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          198:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          199:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          200:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          201:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          202:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          203:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          204:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          205:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          206:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          207:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          208:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          209:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          210:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          211:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          212:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          213:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          214:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          215:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          216:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          217:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          218:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          219:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          220:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          221:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          222:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          223:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          224:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          225:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          226:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          227:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          228:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          229:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          230:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          231:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          232:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          233:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          234:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          235:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          236:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          237:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          238:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          239:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          240:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          241:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          242:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          243:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          244:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          245:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          246:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          247:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          248:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          249:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          250:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          251:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          252:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          253:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          254:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          255:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          256:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          257:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          258:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          259:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          260:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          261:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          262:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          263:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          264:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          265:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          266:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          267:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          268:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          269:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          270:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          271:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          272:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          273:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          274:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          275:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          276:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          277:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          278:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          279:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          280:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          281:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          282:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          283:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          284:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          285:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          286:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          287:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          288:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          289:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          290:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          291:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          292:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          293:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          294:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          295:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          296:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          297:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          298:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          299:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          300:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          301:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          302:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          303:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          304:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          305:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          306:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          307:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          308:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          309:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          310:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          311:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          312:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          313:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          314:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          315:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          316:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          317:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          318:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          319:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          320:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          321:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          322:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          323:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          324:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          325:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          326:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          327:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          328:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          329:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          330:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          331:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          332:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          333:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          334:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          335:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          336:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          337:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          338:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          339:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          340:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          341:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          342:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          343:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          344:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          345:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          346:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          347:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          348:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          349:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          350:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          351:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          352:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          353:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          354:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          355:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          356:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          357:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          358:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          359:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          360:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          361:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          362:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          363:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          364:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          365:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          366:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          367:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          368:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          369:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          370:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          371:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          372:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          373:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          374:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          375:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          376:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          377:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          378:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          379:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          380:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          381:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          382:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          383:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          384:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          385:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          386:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          387:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          388:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          389:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          390:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          391:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          392:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          393:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          394:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          395:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          396:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          397:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          398:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          399:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          400:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          401:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          402:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          403:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          404:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          405:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          406:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          407:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          408:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          409:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          410:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          411:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          412:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          413:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          414:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          415:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          416:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          417:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          418:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          419:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          420:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          421:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          422:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          423:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          424:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          425:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          426:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          427:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          428:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          429:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          430:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          431:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          432:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          433:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          434:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          435:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          436:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          437:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          438:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          439:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          440:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          441:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          442:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          443:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          444:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          445:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          446:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          447:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          448:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          449:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          450:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          451:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          452:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          453:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          454:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          455:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          456:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          457:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          458:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          459:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          460:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          461:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          462:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          463:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          464:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          465:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          466:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          467:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          468:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          469:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          470:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          471:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          472:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          473:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          474:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          475:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          476:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          477:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          478:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          479:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          480:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          481:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          482:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          483:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          484:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          485:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          486:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          487:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          488:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          489:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          490:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          491:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          492:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          493:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          494:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          495:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          496:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          497:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          498:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          499:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          500:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          501:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          502:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          503:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          504:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          505:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          506:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          507:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          508:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          509:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          510:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          511:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          512:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          513:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          514:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          515:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          516:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          517:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          518:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          519:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          520:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          521:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          522:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          523:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          524:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          525:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          526:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          527:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          528:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          529:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          530:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          531:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          532:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          533:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          534:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          535:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          536:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          537:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          538:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          539:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          540:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          541:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          542:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          543:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          544:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          545:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          546:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          547:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          548:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          549:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          550:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          551:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          552:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          553:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          554:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          555:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          556:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          557:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          558:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          559:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          560:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          561:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          562:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          563:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          564:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          565:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          566:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          567:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          568:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          569:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          570:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          571:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          572:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          573:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          574:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          575:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          576:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          577:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          578:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          579:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          580:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          581:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          582:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          583:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          584:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          585:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          586:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          587:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          588:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          589:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          590:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          591:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          592:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          593:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          594:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          595:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          596:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          597:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          598:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          599:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          600:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          601:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          602:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          603:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          604:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          605:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          606:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          607:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          608:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          609:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          610:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          611:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          612:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          613:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          614:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          615:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          616:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          617:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          618:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          619:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          620:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          621:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          622:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          623:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          624:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          625:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          626:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          627:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          628:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          629:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          630:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          631:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          632:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          633:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          634:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          635:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          636:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          637:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          638:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          639:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          640:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          641:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          642:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          643:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          644:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          645:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          646:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          647:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          648:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          649:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          650:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          651:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          652:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          653:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          654:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          655:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          656:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          657:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          658:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          659:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          660:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          661:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          662:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          663:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          664:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          665:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          666:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          667:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          668:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          669:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          670:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          671:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          672:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          673:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          674:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          675:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          676:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          677:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          678:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          679:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          680:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          681:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          682:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          683:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          684:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          685:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          686:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          687:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          688:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          689:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          690:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          691:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          692:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          693:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          694:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          695:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          696:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          697:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          698:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          699:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          700:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          701:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          702:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          703:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          704:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          705:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          706:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          707:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          708:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          709:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          710:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          711:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          712:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          713:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          714:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          715:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          716:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          717:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          718:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          719:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          720:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          721:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          722:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          723:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          724:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          725:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          726:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          727:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          728:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          729:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          730:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          731:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          732:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          733:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          734:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          735:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          736:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          737:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          738:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          739:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          740:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          741:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          742:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          743:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          744:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          745:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          746:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          747:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          748:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          749:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          750:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          751:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          752:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          753:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          754:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          755:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          756:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          757:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          758:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          759:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          760:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          761:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          762:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          763:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          764:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          765:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          766:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          767:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          768:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          769:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          770:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          771:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          772:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          773:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          774:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          775:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          776:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          777:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          778:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          779:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          780:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          781:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          782:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          783:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          784:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          785:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          786:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          787:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          788:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          789:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          790:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          791:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          792:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          793:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          794:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          795:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          796:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          797:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          798:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          799:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          800:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          801:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          802:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          803:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          804:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          805:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          806:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          807:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          808:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          809:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          810:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          811:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          812:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          813:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          814:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          815:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          816:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          817:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          818:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          819:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          820:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          821:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          822:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          823:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          824:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          825:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          826:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          827:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          828:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          829:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          830:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          831:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          832:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          833:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          834:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          835:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          836:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          837:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          838:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          839:
          begin
            cmp[0]<=key_tmp[0];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          840:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          841:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          842:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          843:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          844:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          845:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          846:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          847:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          848:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          849:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          850:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          851:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          852:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          853:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          854:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          855:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          856:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          857:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          858:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          859:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          860:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          861:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          862:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          863:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          864:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          865:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          866:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          867:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          868:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          869:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          870:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          871:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          872:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          873:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          874:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          875:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          876:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          877:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          878:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          879:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          880:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          881:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          882:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          883:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          884:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          885:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          886:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          887:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          888:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          889:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          890:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          891:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          892:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          893:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          894:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          895:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          896:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          897:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          898:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          899:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          900:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          901:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          902:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          903:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          904:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          905:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          906:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          907:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          908:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          909:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          910:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          911:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          912:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          913:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          914:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          915:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          916:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          917:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          918:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          919:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          920:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          921:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          922:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          923:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          924:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          925:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          926:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          927:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          928:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          929:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          930:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          931:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          932:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          933:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          934:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          935:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          936:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          937:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          938:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          939:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          940:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          941:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          942:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          943:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          944:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          945:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          946:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          947:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          948:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          949:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          950:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          951:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          952:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          953:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          954:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          955:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          956:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          957:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          958:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          959:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          960:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          961:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          962:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          963:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          964:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          965:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          966:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          967:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          968:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          969:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          970:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          971:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          972:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          973:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          974:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          975:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          976:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          977:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          978:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          979:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          980:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          981:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          982:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          983:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          984:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          985:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          986:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          987:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          988:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          989:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          990:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          991:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          992:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          993:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          994:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          995:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          996:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          997:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          998:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          999:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1000:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1001:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1002:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1003:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1004:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1005:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1006:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1007:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1008:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1009:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1010:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1011:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1012:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1013:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1014:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1015:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1016:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1017:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1018:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1019:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1020:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1021:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1022:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1023:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1024:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1025:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1026:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1027:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1028:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1029:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1030:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1031:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1032:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1033:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1034:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1035:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1036:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1037:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1038:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1039:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1040:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1041:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1042:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1043:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1044:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1045:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1046:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1047:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1048:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1049:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1050:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1051:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1052:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1053:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1054:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1055:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1056:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1057:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1058:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1059:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1060:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1061:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1062:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1063:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1064:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1065:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1066:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1067:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1068:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1069:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1070:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1071:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1072:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1073:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1074:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1075:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1076:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1077:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1078:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1079:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1080:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1081:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1082:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1083:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1084:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1085:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1086:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1087:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1088:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1089:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1090:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1091:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1092:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1093:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1094:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1095:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1096:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1097:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1098:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1099:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1100:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1101:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1102:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1103:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1104:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1105:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1106:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1107:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1108:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1109:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1110:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1111:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1112:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1113:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1114:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1115:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1116:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1117:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1118:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1119:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1120:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1121:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1122:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1123:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1124:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1125:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1126:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1127:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1128:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1129:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1130:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1131:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1132:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1133:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1134:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1135:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1136:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1137:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1138:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1139:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1140:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1141:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1142:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1143:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1144:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1145:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1146:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1147:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1148:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1149:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1150:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1151:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1152:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1153:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1154:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1155:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1156:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1157:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1158:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1159:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1160:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1161:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1162:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1163:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1164:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1165:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1166:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1167:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1168:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1169:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1170:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1171:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1172:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1173:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1174:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1175:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1176:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1177:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1178:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1179:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1180:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1181:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1182:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1183:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1184:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1185:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1186:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1187:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1188:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1189:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1190:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1191:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1192:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1193:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1194:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1195:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1196:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1197:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1198:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1199:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1200:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1201:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1202:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1203:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1204:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1205:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1206:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1207:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1208:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1209:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1210:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1211:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1212:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1213:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1214:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1215:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1216:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1217:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1218:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1219:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1220:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1221:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1222:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1223:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1224:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1225:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1226:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1227:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1228:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1229:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1230:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1231:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1232:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1233:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1234:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1235:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1236:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1237:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1238:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1239:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1240:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1241:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1242:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1243:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1244:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1245:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1246:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1247:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1248:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1249:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1250:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1251:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1252:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1253:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1254:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1255:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1256:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1257:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1258:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1259:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1260:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1261:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1262:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1263:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1264:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1265:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1266:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1267:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1268:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1269:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1270:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1271:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1272:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1273:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1274:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1275:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1276:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1277:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1278:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1279:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1280:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1281:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1282:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1283:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1284:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1285:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1286:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1287:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1288:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1289:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1290:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1291:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1292:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1293:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1294:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1295:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1296:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1297:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1298:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1299:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1300:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1301:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1302:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1303:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1304:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1305:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1306:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1307:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1308:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1309:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1310:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1311:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1312:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1313:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1314:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1315:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1316:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1317:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1318:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1319:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1320:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1321:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1322:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1323:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1324:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1325:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1326:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1327:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1328:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1329:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1330:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1331:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1332:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1333:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1334:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1335:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1336:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1337:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1338:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1339:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1340:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1341:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1342:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1343:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1344:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1345:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1346:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1347:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1348:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1349:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1350:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1351:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1352:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1353:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1354:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1355:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1356:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1357:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1358:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1359:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1360:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1361:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1362:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1363:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1364:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1365:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1366:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1367:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1368:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1369:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1370:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1371:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1372:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1373:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1374:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1375:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1376:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1377:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1378:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1379:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1380:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1381:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1382:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1383:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1384:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1385:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1386:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1387:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1388:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1389:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1390:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1391:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1392:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1393:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1394:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1395:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1396:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1397:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1398:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1399:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1400:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1401:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1402:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1403:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1404:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1405:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1406:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1407:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1408:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1409:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1410:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1411:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1412:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1413:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1414:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1415:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1416:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1417:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1418:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1419:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1420:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1421:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1422:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1423:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1424:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1425:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1426:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1427:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1428:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1429:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1430:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1431:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1432:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1433:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1434:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1435:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1436:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1437:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1438:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1439:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1440:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1441:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1442:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1443:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1444:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1445:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1446:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1447:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1448:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1449:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1450:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1451:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1452:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1453:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1454:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1455:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1456:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1457:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1458:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1459:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1460:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1461:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1462:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1463:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1464:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1465:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1466:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1467:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1468:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1469:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1470:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1471:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1472:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1473:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1474:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1475:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1476:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1477:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1478:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1479:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1480:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1481:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1482:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1483:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1484:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1485:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1486:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1487:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1488:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1489:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1490:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1491:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1492:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1493:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1494:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1495:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1496:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1497:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1498:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1499:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1500:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1501:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1502:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1503:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1504:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1505:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1506:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1507:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1508:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1509:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1510:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1511:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1512:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1513:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1514:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1515:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1516:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1517:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1518:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1519:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1520:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1521:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1522:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1523:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1524:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1525:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1526:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1527:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          1528:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1529:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1530:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1531:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1532:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1533:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1534:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1535:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1536:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1537:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          1538:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1539:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1540:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1541:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1542:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1543:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1544:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1545:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1546:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1547:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1548:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1549:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1550:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1551:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1552:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1553:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1554:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1555:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1556:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1557:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1558:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1559:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1560:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1561:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1562:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1563:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1564:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1565:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1566:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1567:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1568:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1569:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1570:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1571:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1572:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1573:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1574:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1575:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1576:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1577:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1578:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1579:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1580:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1581:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1582:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1583:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1584:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1585:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1586:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1587:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1588:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1589:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1590:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1591:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1592:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1593:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1594:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1595:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1596:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1597:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1598:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1599:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1600:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1601:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1602:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1603:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1604:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1605:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1606:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1607:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1608:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1609:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1610:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1611:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1612:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1613:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1614:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1615:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1616:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1617:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1618:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1619:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1620:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1621:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1622:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1623:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1624:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1625:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1626:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1627:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1628:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1629:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1630:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1631:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1632:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1633:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1634:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1635:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1636:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1637:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1638:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1639:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1640:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1641:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1642:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1643:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1644:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1645:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1646:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1647:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          1648:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1649:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1650:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1651:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1652:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1653:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1654:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1655:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1656:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1657:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          1658:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1659:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1660:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          1661:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1662:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1663:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1664:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          1665:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          1666:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          1667:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          1668:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1669:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          1670:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1671:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1672:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1673:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          1674:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1675:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1676:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1677:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          1678:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1679:
          begin
            cmp[0]<=key_tmp[1];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1680:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1681:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1682:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1683:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1684:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1685:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1686:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1687:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1688:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1689:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1690:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1691:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1692:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1693:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1694:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1695:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1696:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1697:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1698:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1699:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1700:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          1701:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          1702:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1703:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1704:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          1705:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1706:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1707:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1708:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          1709:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1710:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1711:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1712:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1713:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1714:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1715:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1716:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1717:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1718:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1719:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1720:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          1721:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          1722:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1723:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1724:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          1725:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1726:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1727:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1728:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          1729:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1730:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1731:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1732:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1733:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1734:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1735:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1736:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1737:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1738:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1739:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1740:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          1741:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          1742:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1743:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1744:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          1745:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1746:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1747:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1748:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          1749:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1750:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1751:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1752:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1753:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1754:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1755:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1756:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1757:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1758:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1759:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1760:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          1761:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          1762:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          1763:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1764:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          1765:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1766:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1767:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1768:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          1769:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1770:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1771:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1772:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          1773:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1774:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1775:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1776:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1777:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1778:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1779:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1780:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          1781:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          1782:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          1783:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1784:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          1785:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1786:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1787:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1788:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          1789:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1790:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1791:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1792:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          1793:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1794:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1795:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1796:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1797:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1798:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1799:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1800:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1801:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1802:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1803:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1804:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1805:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1806:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1807:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1808:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1809:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1810:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1811:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1812:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1813:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1814:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1815:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1816:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1817:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1818:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1819:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1820:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1821:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1822:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1823:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1824:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1825:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1826:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1827:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1828:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1829:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1830:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1831:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1832:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1833:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1834:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1835:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1836:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1837:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1838:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1839:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1840:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1841:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1842:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1843:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1844:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1845:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1846:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1847:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1848:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1849:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1850:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1851:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1852:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1853:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1854:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1855:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1856:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1857:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1858:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1859:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1860:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1861:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1862:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1863:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1864:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1865:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1866:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1867:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1868:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1869:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1870:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1871:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1872:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1873:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1874:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1875:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1876:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1877:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1878:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1879:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1880:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1881:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1882:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1883:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1884:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1885:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1886:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1887:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          1888:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1889:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1890:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1891:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1892:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1893:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1894:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1895:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1896:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1897:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          1898:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1899:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1900:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          1901:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1902:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1903:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1904:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          1905:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          1906:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          1907:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          1908:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1909:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          1910:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1911:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1912:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1913:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          1914:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1915:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1916:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1917:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          1918:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1919:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1920:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          1921:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          1922:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1923:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1924:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          1925:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1926:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1927:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1928:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          1929:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1930:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1931:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1932:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1933:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1934:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1935:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1936:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1937:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1938:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1939:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1940:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1941:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1942:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1943:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1944:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1945:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          1946:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1947:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1948:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1949:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          1950:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1951:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1952:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1953:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1954:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1955:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1956:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1957:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1958:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1959:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1960:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          1961:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          1962:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1963:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1964:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          1965:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          1966:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1967:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1968:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          1969:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          1970:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          1971:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          1972:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1973:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1974:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          1975:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1976:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1977:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1978:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          1979:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          1980:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          1981:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          1982:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          1983:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          1984:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          1985:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          1986:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          1987:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          1988:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          1989:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          1990:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          1991:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          1992:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          1993:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          1994:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          1995:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          1996:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          1997:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          1998:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          1999:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2000:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2001:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2002:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2003:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2004:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2005:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2006:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2007:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2008:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2009:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2010:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2011:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2012:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2013:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2014:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2015:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2016:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2017:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2018:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2019:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2020:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2021:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2022:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2023:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2024:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2025:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2026:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2027:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2028:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2029:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2030:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2031:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2032:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2033:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2034:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2035:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2036:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2037:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2038:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2039:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2040:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2041:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2042:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2043:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2044:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2045:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2046:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2047:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2048:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2049:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2050:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2051:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2052:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2053:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2054:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2055:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2056:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2057:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2058:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2059:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2060:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2061:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2062:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2063:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2064:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2065:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2066:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2067:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2068:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2069:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2070:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2071:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2072:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2073:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2074:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2075:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2076:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2077:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2078:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2079:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2080:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2081:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2082:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2083:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2084:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2085:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2086:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2087:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2088:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2089:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2090:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2091:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2092:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2093:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2094:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2095:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2096:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2097:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2098:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2099:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2100:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2101:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2102:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2103:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2104:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2105:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2106:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2107:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2108:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2109:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2110:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2111:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2112:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2113:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2114:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2115:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2116:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2117:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2118:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2119:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2120:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2121:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2122:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2123:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2124:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2125:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2126:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2127:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2128:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2129:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2130:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2131:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2132:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2133:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2134:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2135:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2136:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2137:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2138:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2139:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2140:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2141:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2142:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2143:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2144:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2145:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2146:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2147:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2148:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2149:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2150:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2151:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2152:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2153:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2154:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2155:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2156:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2157:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2158:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2159:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2160:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2161:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2162:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2163:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2164:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2165:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2166:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2167:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2168:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2169:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2170:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2171:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2172:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2173:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2174:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2175:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2176:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2177:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2178:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2179:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2180:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2181:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2182:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2183:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2184:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2185:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2186:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2187:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2188:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2189:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2190:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2191:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2192:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2193:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2194:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2195:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2196:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2197:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2198:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2199:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2200:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2201:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2202:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2203:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2204:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2205:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2206:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2207:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2208:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2209:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2210:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2211:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2212:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2213:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2214:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2215:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2216:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2217:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2218:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2219:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2220:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2221:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2222:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2223:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2224:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2225:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2226:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2227:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2228:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2229:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2230:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2231:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2232:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2233:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2234:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2235:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2236:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2237:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2238:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2239:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2240:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2241:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2242:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2243:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2244:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2245:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2246:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2247:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2248:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2249:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2250:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2251:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2252:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2253:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2254:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2255:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2256:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2257:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2258:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2259:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2260:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2261:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2262:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2263:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2264:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2265:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2266:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2267:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2268:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2269:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2270:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2271:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2272:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2273:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2274:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2275:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2276:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2277:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2278:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2279:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2280:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2281:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2282:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2283:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2284:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2285:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2286:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2287:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2288:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2289:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2290:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2291:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2292:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2293:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2294:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2295:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2296:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2297:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2298:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2299:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2300:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2301:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2302:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2303:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2304:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2305:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2306:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2307:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2308:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2309:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2310:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2311:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2312:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2313:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2314:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2315:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2316:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2317:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2318:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2319:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2320:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2321:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2322:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2323:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2324:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2325:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2326:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2327:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2328:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2329:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2330:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2331:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2332:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2333:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2334:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2335:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2336:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2337:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2338:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2339:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2340:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2341:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2342:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2343:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2344:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2345:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2346:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2347:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2348:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2349:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2350:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2351:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2352:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2353:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2354:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2355:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2356:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2357:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2358:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2359:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2360:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2361:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2362:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2363:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2364:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2365:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2366:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2367:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2368:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2369:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2370:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2371:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          2372:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2373:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2374:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2375:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2376:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2377:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2378:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          2379:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2380:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2381:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2382:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2383:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2384:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2385:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2386:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2387:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2388:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2389:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2390:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2391:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2392:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2393:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2394:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2395:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2396:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2397:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2398:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2399:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2400:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2401:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2402:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2403:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2404:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2405:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2406:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2407:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2408:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2409:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2410:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2411:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2412:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2413:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2414:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2415:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2416:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2417:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2418:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2419:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2420:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2421:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2422:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2423:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2424:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2425:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2426:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2427:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2428:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2429:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2430:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2431:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2432:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2433:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2434:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2435:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2436:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2437:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2438:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2439:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2440:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2441:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2442:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2443:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2444:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2445:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2446:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2447:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2448:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2449:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2450:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2451:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2452:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2453:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2454:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2455:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2456:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2457:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2458:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2459:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2460:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2461:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2462:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2463:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2464:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2465:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2466:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2467:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2468:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2469:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2470:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2471:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2472:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2473:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2474:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2475:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2476:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2477:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2478:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2479:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2480:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2481:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2482:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2483:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2484:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2485:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2486:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2487:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2488:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2489:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2490:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2491:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          2492:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2493:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2494:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2495:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2496:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2497:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2498:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          2499:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2500:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2501:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          2502:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2503:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2504:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2505:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          2506:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2507:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2508:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          2509:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          2510:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          2511:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          2512:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2513:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2514:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          2515:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2516:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2517:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2518:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          2519:
          begin
            cmp[0]<=key_tmp[2];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2520:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2521:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2522:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2523:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2524:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2525:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2526:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2527:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2528:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2529:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2530:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2531:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2532:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2533:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2534:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2535:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2536:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2537:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2538:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2539:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2540:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2541:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2542:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2543:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2544:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2545:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2546:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2547:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2548:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2549:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2550:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2551:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2552:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2553:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2554:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2555:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2556:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2557:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2558:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2559:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2560:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2561:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2562:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2563:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2564:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2565:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2566:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2567:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2568:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2569:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2570:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2571:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2572:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2573:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2574:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2575:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2576:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2577:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2578:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2579:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2580:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2581:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2582:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2583:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2584:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2585:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2586:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2587:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2588:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2589:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2590:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2591:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2592:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2593:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2594:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2595:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2596:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2597:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2598:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2599:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2600:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2601:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2602:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2603:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2604:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2605:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2606:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2607:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2608:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2609:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2610:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2611:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2612:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2613:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2614:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2615:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2616:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2617:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2618:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2619:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2620:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2621:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2622:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2623:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2624:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2625:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2626:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2627:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2628:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2629:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2630:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2631:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2632:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2633:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2634:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2635:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2636:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2637:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2638:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2639:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2640:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2641:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2642:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2643:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2644:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2645:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2646:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2647:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2648:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2649:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2650:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2651:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2652:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2653:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2654:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2655:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2656:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2657:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2658:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2659:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2660:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2661:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2662:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2663:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2664:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2665:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2666:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2667:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2668:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2669:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2670:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2671:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2672:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2673:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2674:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2675:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2676:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2677:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2678:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2679:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2680:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2681:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2682:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2683:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2684:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2685:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2686:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2687:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2688:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2689:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2690:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2691:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2692:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2693:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2694:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2695:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2696:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2697:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2698:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2699:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2700:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2701:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2702:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2703:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2704:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2705:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2706:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2707:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2708:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2709:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2710:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2711:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2712:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2713:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2714:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2715:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2716:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2717:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2718:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2719:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2720:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2721:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2722:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2723:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2724:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2725:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2726:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2727:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2728:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2729:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2730:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2731:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2732:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2733:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2734:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2735:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2736:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2737:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2738:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2739:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2740:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2741:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2742:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2743:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2744:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2745:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          2746:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2747:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2748:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2749:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          2750:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2751:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2752:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2753:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2754:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2755:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2756:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2757:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2758:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2759:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2760:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2761:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2762:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2763:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2764:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2765:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2766:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2767:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2768:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2769:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2770:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2771:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2772:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2773:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2774:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2775:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2776:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2777:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2778:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2779:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2780:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2781:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2782:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2783:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2784:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2785:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2786:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2787:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2788:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2789:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2790:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2791:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2792:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2793:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2794:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2795:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2796:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2797:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2798:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2799:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2800:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2801:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2802:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2803:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2804:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2805:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2806:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2807:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2808:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2809:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2810:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2811:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2812:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2813:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2814:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2815:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2816:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2817:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2818:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2819:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2820:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2821:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2822:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2823:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2824:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2825:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2826:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2827:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2828:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2829:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2830:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2831:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2832:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2833:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2834:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2835:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2836:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2837:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2838:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2839:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2840:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2841:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2842:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2843:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2844:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2845:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2846:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2847:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2848:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2849:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2850:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2851:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          2852:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2853:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2854:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2855:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2856:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2857:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2858:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          2859:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2860:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2861:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          2862:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2863:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2864:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2865:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          2866:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2867:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2868:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          2869:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          2870:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          2871:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          2872:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2873:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2874:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          2875:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2876:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2877:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2878:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          2879:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2880:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2881:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2882:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2883:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2884:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2885:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2886:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2887:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2888:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2889:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2890:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2891:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2892:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2893:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2894:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2895:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2896:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2897:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2898:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2899:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2900:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2901:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2902:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2903:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2904:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2905:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2906:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2907:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2908:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2909:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2910:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2911:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2912:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2913:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2914:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2915:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2916:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2917:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2918:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2919:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2920:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2921:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2922:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2923:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2924:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2925:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2926:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2927:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2928:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2929:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2930:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2931:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2932:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2933:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2934:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          2935:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2936:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2937:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2938:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2939:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2940:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2941:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2942:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2943:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2944:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2945:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2946:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2947:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2948:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2949:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2950:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2951:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2952:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2953:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2954:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2955:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          2956:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2957:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2958:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2959:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          2960:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2961:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2962:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2963:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          2964:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2965:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2966:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2967:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          2968:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2969:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2970:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2971:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          2972:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2973:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2974:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2975:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          2976:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          2977:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          2978:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          2979:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          2980:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          2981:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          2982:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          2983:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          2984:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          2985:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          2986:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          2987:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          2988:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          2989:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          2990:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          2991:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          2992:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          2993:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          2994:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          2995:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          2996:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          2997:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          2998:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          2999:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3000:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3001:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3002:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3003:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3004:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3005:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3006:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3007:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3008:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3009:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3010:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3011:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3012:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3013:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3014:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3015:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3016:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3017:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3018:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3019:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3020:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3021:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3022:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3023:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3024:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3025:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3026:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3027:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3028:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3029:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3030:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3031:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3032:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3033:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3034:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3035:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3036:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3037:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3038:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3039:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3040:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3041:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3042:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3043:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3044:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3045:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3046:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3047:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3048:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3049:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3050:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3051:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3052:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3053:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3054:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3055:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3056:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3057:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3058:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3059:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3060:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3061:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3062:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3063:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3064:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3065:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3066:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3067:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3068:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3069:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3070:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3071:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3072:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3073:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3074:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3075:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3076:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3077:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3078:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3079:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3080:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3081:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3082:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3083:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3084:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3085:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3086:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3087:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3088:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3089:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3090:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3091:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3092:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3093:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3094:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3095:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3096:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3097:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3098:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3099:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3100:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3101:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3102:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3103:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3104:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3105:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3106:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3107:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3108:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3109:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3110:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3111:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3112:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3113:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3114:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3115:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3116:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3117:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3118:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3119:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3120:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3121:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3122:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3123:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3124:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3125:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3126:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3127:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3128:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3129:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3130:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3131:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3132:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3133:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3134:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3135:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3136:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3137:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3138:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3139:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3140:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3141:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3142:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3143:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3144:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3145:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3146:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3147:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3148:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3149:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3150:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3151:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3152:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3153:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3154:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3155:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3156:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3157:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3158:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3159:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3160:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3161:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3162:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3163:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3164:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3165:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3166:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3167:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3168:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3169:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3170:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3171:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3172:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3173:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3174:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3175:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3176:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3177:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3178:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3179:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3180:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3181:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3182:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3183:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3184:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3185:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3186:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3187:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3188:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3189:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3190:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3191:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3192:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3193:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3194:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3195:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3196:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3197:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3198:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3199:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3200:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3201:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3202:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3203:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3204:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3205:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3206:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3207:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3208:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3209:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3210:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3211:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3212:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3213:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3214:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3215:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          3216:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3217:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3218:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3219:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          3220:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3221:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3222:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3223:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3224:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3225:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3226:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3227:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3228:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3229:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3230:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3231:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3232:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3233:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3234:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3235:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3236:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3237:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3238:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3239:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3240:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3241:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3242:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3243:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3244:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3245:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3246:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3247:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3248:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3249:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3250:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3251:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3252:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3253:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3254:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3255:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3256:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3257:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3258:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3259:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3260:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3261:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3262:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3263:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3264:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3265:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3266:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3267:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3268:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3269:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3270:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3271:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3272:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3273:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3274:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3275:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3276:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3277:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3278:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3279:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3280:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3281:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3282:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3283:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3284:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3285:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3286:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3287:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3288:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3289:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3290:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3291:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3292:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3293:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3294:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3295:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3296:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3297:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3298:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3299:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3300:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3301:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3302:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3303:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3304:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3305:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3306:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3307:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3308:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3309:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3310:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3311:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3312:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3313:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3314:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3315:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3316:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3317:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3318:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3319:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3320:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3321:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3322:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3323:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3324:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3325:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3326:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3327:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3328:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3329:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3330:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3331:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3332:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3333:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3334:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3335:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          3336:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3337:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3338:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3339:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          3340:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3341:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3342:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          3343:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3344:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3345:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3346:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          3347:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3348:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3349:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3350:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          3351:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3352:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          3353:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          3354:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          3355:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          3356:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3357:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3358:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3359:
          begin
            cmp[0]<=key_tmp[3];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          3360:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3361:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3362:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3363:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3364:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3365:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3366:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3367:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3368:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3369:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3370:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3371:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3372:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3373:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3374:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3375:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3376:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3377:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3378:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3379:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3380:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3381:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3382:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3383:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3384:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3385:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3386:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3387:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3388:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3389:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3390:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3391:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3392:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3393:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3394:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3395:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3396:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3397:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3398:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3399:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3400:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3401:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3402:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3403:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3404:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3405:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3406:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3407:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3408:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3409:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3410:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3411:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3412:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3413:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3414:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3415:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3416:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3417:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3418:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3419:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3420:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3421:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3422:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3423:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3424:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3425:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3426:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3427:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3428:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3429:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3430:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3431:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3432:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3433:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3434:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3435:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3436:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3437:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3438:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3439:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3440:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3441:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3442:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3443:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3444:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3445:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3446:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3447:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3448:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3449:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3450:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3451:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3452:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3453:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3454:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3455:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3456:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3457:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3458:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3459:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3460:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3461:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3462:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3463:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3464:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3465:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3466:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3467:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3468:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3469:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3470:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3471:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3472:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3473:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3474:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3475:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3476:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3477:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3478:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3479:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3480:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3481:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3482:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3483:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3484:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3485:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3486:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3487:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3488:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3489:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3490:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3491:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3492:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3493:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3494:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3495:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3496:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3497:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3498:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3499:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3500:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3501:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3502:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3503:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3504:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3505:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3506:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3507:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3508:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3509:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3510:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3511:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3512:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3513:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3514:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3515:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3516:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3517:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3518:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3519:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3520:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3521:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3522:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3523:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3524:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3525:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3526:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3527:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3528:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3529:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3530:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3531:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3532:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3533:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3534:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3535:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3536:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3537:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3538:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3539:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3540:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3541:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3542:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3543:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3544:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3545:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3546:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3547:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3548:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3549:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3550:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3551:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3552:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3553:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3554:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3555:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3556:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3557:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3558:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3559:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3560:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3561:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3562:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3563:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3564:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3565:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3566:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3567:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3568:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3569:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3570:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3571:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3572:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3573:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3574:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3575:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3576:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3577:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3578:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3579:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3580:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3581:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3582:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3583:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3584:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3585:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3586:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3587:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3588:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3589:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3590:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3591:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3592:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3593:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3594:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3595:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3596:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3597:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3598:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3599:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3600:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3601:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3602:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3603:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3604:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3605:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3606:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3607:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3608:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3609:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3610:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3611:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3612:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3613:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3614:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3615:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3616:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3617:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3618:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3619:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3620:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3621:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3622:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3623:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3624:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3625:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3626:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3627:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3628:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3629:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3630:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3631:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3632:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3633:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3634:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3635:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3636:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3637:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3638:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3639:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3640:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3641:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3642:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3643:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3644:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3645:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3646:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3647:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3648:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3649:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3650:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3651:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3652:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3653:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3654:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3655:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3656:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3657:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3658:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3659:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3660:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3661:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3662:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3663:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3664:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3665:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3666:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3667:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3668:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3669:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3670:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3671:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3672:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3673:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3674:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3675:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3676:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3677:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3678:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3679:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3680:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3681:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3682:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3683:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3684:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3685:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3686:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3687:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3688:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3689:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3690:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3691:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3692:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3693:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3694:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3695:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3696:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3697:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3698:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3699:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3700:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3701:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3702:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3703:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3704:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3705:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3706:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3707:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3708:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3709:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3710:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3711:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3712:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3713:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3714:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3715:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3716:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3717:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3718:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3719:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3720:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3721:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3722:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3723:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3724:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3725:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3726:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3727:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3728:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3729:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3730:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3731:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3732:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3733:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3734:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3735:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3736:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3737:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3738:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3739:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3740:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3741:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3742:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3743:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3744:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3745:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3746:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3747:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3748:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3749:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3750:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3751:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3752:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3753:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3754:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3755:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3756:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3757:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3758:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3759:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3760:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3761:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3762:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3763:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3764:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3765:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3766:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3767:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3768:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3769:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3770:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3771:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3772:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3773:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3774:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3775:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3776:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3777:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3778:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3779:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3780:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3781:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3782:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3783:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3784:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3785:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3786:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3787:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3788:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3789:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3790:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3791:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3792:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3793:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3794:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3795:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3796:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3797:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3798:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3799:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3800:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3801:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3802:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3803:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3804:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3805:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3806:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3807:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3808:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3809:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3810:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3811:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3812:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3813:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3814:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3815:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3816:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3817:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3818:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3819:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3820:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3821:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3822:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3823:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3824:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3825:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3826:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3827:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3828:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3829:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3830:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3831:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3832:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3833:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3834:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3835:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          3836:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3837:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3838:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3839:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          3840:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3841:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3842:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3843:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3844:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3845:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3846:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3847:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3848:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3849:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3850:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3851:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3852:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3853:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3854:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3855:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3856:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3857:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3858:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3859:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3860:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3861:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3862:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3863:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3864:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3865:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3866:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3867:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3868:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3869:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3870:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3871:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3872:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3873:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3874:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3875:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3876:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3877:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3878:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3879:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3880:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3881:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3882:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3883:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3884:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3885:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3886:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3887:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3888:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3889:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3890:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3891:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3892:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3893:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3894:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3895:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3896:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3897:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3898:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3899:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3900:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3901:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3902:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3903:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3904:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3905:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3906:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3907:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3908:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3909:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3910:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3911:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3912:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3913:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3914:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3915:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          3916:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3917:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3918:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3919:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          3920:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3921:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3922:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3923:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3924:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3925:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3926:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3927:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3928:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3929:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3930:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3931:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3932:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3933:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3934:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3935:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3936:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3937:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3938:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3939:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3940:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          3941:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3942:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3943:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          3944:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          3945:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3946:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3947:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          3948:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3949:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3950:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3951:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          3952:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3953:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3954:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3955:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          3956:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          3957:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          3958:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          3959:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          3960:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          3961:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          3962:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          3963:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          3964:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          3965:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3966:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3967:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3968:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          3969:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3970:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3971:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3972:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          3973:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3974:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3975:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3976:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          3977:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3978:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3979:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          3980:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          3981:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          3982:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          3983:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          3984:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          3985:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          3986:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          3987:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          3988:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          3989:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          3990:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          3991:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          3992:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          3993:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          3994:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          3995:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          3996:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          3997:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          3998:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          3999:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          4000:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4001:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4002:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4003:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4004:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4005:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4006:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4007:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4008:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4009:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4010:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          4011:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4012:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4013:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4014:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          4015:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          4016:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4017:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4018:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4019:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          4020:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4021:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4022:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4023:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4024:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4025:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4026:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4027:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4028:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4029:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4030:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          4031:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4032:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4033:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4034:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          4035:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          4036:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4037:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4038:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4039:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          4040:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4041:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4042:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4043:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4044:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4045:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4046:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4047:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4048:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4049:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4050:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4051:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4052:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4053:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4054:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4055:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4056:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4057:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4058:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4059:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4060:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4061:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4062:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4063:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4064:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4065:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4066:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4067:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4068:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4069:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4070:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4071:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          4072:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4073:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4074:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4075:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          4076:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4077:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4078:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          4079:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          4080:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4081:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4082:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4083:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4084:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4085:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4086:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          4087:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4088:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4089:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4090:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          4091:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4092:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4093:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          4094:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          4095:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          4096:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4097:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4098:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4099:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          4100:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4101:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4102:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4103:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4104:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4105:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4106:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          4107:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4108:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4109:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4110:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          4111:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4112:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4113:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          4114:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          4115:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          4116:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4117:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4118:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4119:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          4120:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4121:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4122:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4123:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4124:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4125:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4126:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4127:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4128:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4129:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4130:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          4131:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4132:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4133:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4134:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          4135:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          4136:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4137:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4138:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4139:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          4140:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4141:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4142:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4143:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4144:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4145:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4146:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4147:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4148:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4149:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4150:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          4151:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4152:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4153:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4154:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          4155:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          4156:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4157:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4158:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4159:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          4160:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4161:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4162:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4163:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4164:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4165:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4166:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4167:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4168:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4169:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4170:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4171:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4172:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4173:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4174:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4175:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4176:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4177:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4178:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4179:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4180:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4181:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4182:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4183:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          4184:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4185:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4186:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4187:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          4188:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4189:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4190:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4191:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          4192:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4193:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4194:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4195:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          4196:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          4197:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          4198:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          4199:
          begin
            cmp[0]<=key_tmp[4];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          4200:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4201:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4202:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4203:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4204:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4205:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4206:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4207:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4208:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4209:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4210:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4211:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4212:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4213:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4214:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4215:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4216:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4217:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4218:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4219:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4220:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4221:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4222:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4223:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4224:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4225:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4226:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4227:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4228:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4229:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4230:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4231:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4232:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4233:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4234:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4235:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4236:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4237:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4238:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4239:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4240:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4241:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4242:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4243:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4244:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4245:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4246:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4247:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4248:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4249:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4250:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4251:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4252:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4253:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4254:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4255:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4256:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4257:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4258:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4259:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4260:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4261:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4262:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4263:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4264:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4265:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4266:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4267:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4268:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4269:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4270:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4271:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4272:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4273:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4274:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4275:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4276:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4277:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4278:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4279:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4280:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4281:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4282:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4283:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4284:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4285:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4286:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4287:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4288:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4289:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4290:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4291:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4292:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4293:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4294:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4295:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4296:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4297:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4298:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4299:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4300:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4301:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4302:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4303:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4304:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4305:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4306:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4307:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4308:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4309:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4310:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4311:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4312:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4313:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4314:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4315:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4316:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4317:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4318:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4319:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4320:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4321:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4322:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4323:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4324:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4325:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4326:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4327:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4328:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4329:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4330:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4331:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4332:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4333:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4334:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4335:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4336:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4337:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4338:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4339:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4340:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4341:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4342:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4343:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4344:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4345:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4346:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4347:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4348:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4349:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4350:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4351:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4352:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4353:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4354:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4355:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4356:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4357:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4358:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4359:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4360:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4361:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4362:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4363:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4364:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4365:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4366:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4367:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4368:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4369:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4370:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4371:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4372:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4373:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4374:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4375:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4376:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4377:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4378:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4379:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4380:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4381:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4382:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4383:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4384:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4385:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4386:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4387:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4388:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4389:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4390:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4391:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4392:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4393:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4394:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4395:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4396:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4397:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4398:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4399:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4400:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4401:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4402:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4403:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4404:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4405:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4406:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4407:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4408:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4409:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4410:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4411:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4412:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4413:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4414:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4415:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4416:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4417:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4418:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4419:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4420:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4421:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4422:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4423:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4424:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4425:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4426:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4427:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4428:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4429:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4430:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4431:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4432:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4433:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4434:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4435:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4436:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4437:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4438:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4439:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4440:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4441:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4442:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4443:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4444:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4445:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4446:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4447:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4448:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4449:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4450:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4451:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4452:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4453:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4454:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4455:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4456:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4457:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4458:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4459:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4460:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4461:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4462:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4463:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4464:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4465:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4466:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4467:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4468:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4469:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4470:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4471:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4472:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4473:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4474:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4475:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4476:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4477:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4478:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4479:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4480:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4481:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4482:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4483:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4484:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4485:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4486:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4487:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4488:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4489:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4490:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4491:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4492:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4493:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4494:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4495:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4496:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4497:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4498:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4499:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4500:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4501:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4502:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4503:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4504:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4505:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4506:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4507:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4508:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4509:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4510:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4511:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4512:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4513:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4514:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4515:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4516:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4517:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4518:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4519:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4520:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4521:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4522:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4523:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4524:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4525:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4526:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4527:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4528:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4529:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4530:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4531:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4532:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4533:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4534:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4535:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4536:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4537:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4538:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4539:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4540:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4541:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4542:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4543:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4544:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4545:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4546:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4547:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4548:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4549:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4550:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4551:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4552:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4553:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4554:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4555:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4556:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4557:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4558:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4559:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4560:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4561:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4562:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4563:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4564:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4565:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4566:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4567:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4568:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4569:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4570:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4571:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4572:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4573:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4574:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4575:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4576:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4577:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4578:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4579:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4580:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4581:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4582:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4583:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4584:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4585:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4586:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4587:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4588:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4589:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4590:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4591:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4592:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4593:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4594:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4595:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4596:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4597:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4598:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4599:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4600:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4601:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4602:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4603:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4604:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4605:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4606:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4607:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4608:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4609:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4610:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4611:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4612:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4613:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4614:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4615:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4616:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4617:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4618:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4619:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4620:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4621:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4622:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4623:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4624:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4625:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4626:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4627:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4628:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4629:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4630:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4631:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4632:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4633:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4634:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4635:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4636:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4637:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4638:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4639:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4640:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4641:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4642:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4643:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4644:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4645:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4646:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4647:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4648:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4649:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4650:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4651:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4652:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4653:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4654:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4655:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4656:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4657:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4658:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4659:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4660:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4661:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4662:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4663:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4664:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4665:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4666:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4667:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4668:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4669:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4670:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4671:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4672:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4673:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4674:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4675:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4676:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4677:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4678:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4679:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4680:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4681:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4682:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4683:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4684:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4685:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4686:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4687:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4688:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4689:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4690:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4691:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4692:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4693:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4694:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4695:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4696:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4697:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4698:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4699:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4700:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4701:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4702:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4703:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4704:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4705:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4706:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4707:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4708:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4709:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4710:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4711:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4712:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4713:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4714:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4715:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4716:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4717:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4718:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4719:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4720:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4721:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4722:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4723:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4724:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4725:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4726:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4727:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4728:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4729:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4730:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4731:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4732:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4733:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4734:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4735:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4736:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4737:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4738:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4739:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4740:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4741:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4742:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4743:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4744:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4745:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4746:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4747:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4748:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4749:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4750:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4751:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4752:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4753:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4754:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4755:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[7];
          end
          4756:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4757:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4758:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4759:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[6];
          end
          4760:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4761:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4762:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4763:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4764:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4765:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4766:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4767:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4768:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4769:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4770:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4771:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4772:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4773:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4774:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4775:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4776:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4777:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4778:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4779:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4780:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4781:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4782:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4783:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4784:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4785:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4786:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4787:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4788:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4789:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4790:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4791:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4792:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4793:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4794:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4795:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4796:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4797:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4798:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4799:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4800:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4801:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4802:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4803:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4804:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4805:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4806:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4807:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4808:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4809:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4810:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4811:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4812:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4813:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4814:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4815:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4816:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4817:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4818:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4819:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4820:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4821:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4822:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4823:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4824:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4825:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4826:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4827:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4828:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4829:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4830:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4831:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4832:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4833:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4834:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4835:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4836:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4837:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4838:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4839:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4840:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4841:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4842:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4843:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4844:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4845:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4846:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4847:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4848:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4849:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4850:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4851:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4852:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4853:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4854:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4855:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4856:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4857:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4858:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4859:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4860:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4861:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4862:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4863:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4864:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4865:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4866:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4867:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4868:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4869:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4870:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4871:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4872:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4873:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4874:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4875:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          4876:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4877:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4878:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4879:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          4880:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4881:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4882:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4883:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          4884:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4885:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4886:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4887:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          4888:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4889:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4890:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4891:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          4892:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4893:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4894:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4895:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          4896:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          4897:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          4898:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          4899:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          4900:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4901:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4902:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4903:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4904:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4905:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4906:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4907:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4908:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4909:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4910:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4911:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4912:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4913:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4914:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4915:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4916:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4917:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4918:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4919:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4920:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4921:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4922:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4923:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4924:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4925:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4926:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4927:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4928:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4929:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4930:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4931:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4932:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4933:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4934:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4935:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4936:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4937:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4938:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4939:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4940:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4941:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4942:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4943:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4944:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4945:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          4946:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4947:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4948:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4949:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          4950:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4951:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4952:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4953:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4954:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4955:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4956:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4957:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4958:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4959:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4960:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4961:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          4962:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4963:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4964:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4965:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          4966:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4967:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4968:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          4969:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          4970:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          4971:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          4972:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4973:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4974:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          4975:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4976:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4977:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4978:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          4979:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          4980:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          4981:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          4982:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          4983:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          4984:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          4985:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          4986:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          4987:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          4988:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          4989:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          4990:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          4991:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          4992:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          4993:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          4994:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          4995:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          4996:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          4997:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          4998:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          4999:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          5000:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5001:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5002:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5003:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          5004:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5005:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5006:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5007:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          5008:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5009:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5010:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5011:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          5012:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5013:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5014:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5015:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          5016:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          5017:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          5018:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          5019:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          5020:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5021:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5022:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5023:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5024:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5025:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5026:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5027:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5028:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5029:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5030:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5031:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5032:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5033:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5034:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5035:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5036:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5037:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5038:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5039:
          begin
            cmp[0]<=key_tmp[5];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5040:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5041:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5042:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5043:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5044:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5045:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5046:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5047:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5048:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5049:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5050:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5051:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5052:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5053:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5054:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5055:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5056:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5057:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5058:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5059:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5060:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5061:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5062:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5063:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5064:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5065:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5066:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5067:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5068:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5069:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5070:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5071:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5072:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5073:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5074:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5075:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5076:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5077:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5078:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5079:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5080:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5081:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5082:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5083:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5084:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5085:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5086:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5087:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5088:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5089:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5090:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5091:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5092:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5093:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5094:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5095:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5096:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5097:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5098:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5099:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5100:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5101:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5102:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5103:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5104:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5105:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5106:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5107:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5108:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5109:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5110:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5111:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5112:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5113:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5114:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5115:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5116:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5117:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5118:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5119:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5120:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5121:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5122:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5123:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5124:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5125:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5126:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5127:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5128:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5129:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5130:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5131:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5132:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5133:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5134:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5135:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5136:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5137:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5138:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5139:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5140:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5141:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5142:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5143:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5144:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5145:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5146:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5147:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5148:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5149:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5150:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5151:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5152:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5153:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5154:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5155:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5156:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5157:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5158:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5159:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5160:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5161:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5162:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5163:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5164:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5165:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5166:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5167:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5168:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5169:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5170:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5171:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5172:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5173:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5174:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5175:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5176:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5177:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5178:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5179:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5180:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5181:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5182:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5183:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5184:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5185:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5186:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5187:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5188:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5189:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5190:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5191:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5192:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5193:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5194:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5195:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5196:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5197:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5198:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5199:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5200:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5201:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5202:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5203:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5204:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5205:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5206:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5207:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5208:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5209:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5210:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5211:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5212:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5213:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5214:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5215:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5216:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5217:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5218:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5219:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5220:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5221:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5222:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5223:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5224:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5225:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5226:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5227:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5228:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5229:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5230:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5231:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5232:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5233:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5234:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5235:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5236:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5237:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5238:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5239:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5240:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5241:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5242:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5243:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5244:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5245:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5246:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5247:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5248:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5249:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5250:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5251:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5252:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5253:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5254:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5255:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5256:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5257:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5258:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5259:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5260:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5261:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5262:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5263:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5264:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5265:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5266:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5267:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5268:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5269:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5270:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5271:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5272:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5273:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5274:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5275:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5276:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5277:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5278:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5279:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5280:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5281:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5282:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5283:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5284:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5285:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5286:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5287:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5288:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5289:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5290:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5291:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5292:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5293:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5294:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5295:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5296:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5297:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5298:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5299:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5300:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5301:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5302:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5303:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5304:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5305:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5306:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5307:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5308:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5309:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5310:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5311:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5312:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5313:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5314:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5315:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5316:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5317:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5318:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5319:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5320:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5321:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5322:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5323:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5324:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5325:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5326:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5327:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5328:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5329:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5330:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5331:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5332:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5333:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5334:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5335:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5336:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5337:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5338:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5339:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5340:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5341:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5342:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5343:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5344:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5345:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5346:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5347:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5348:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5349:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5350:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5351:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5352:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5353:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5354:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5355:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5356:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5357:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5358:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5359:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5360:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5361:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5362:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5363:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5364:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5365:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5366:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5367:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5368:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5369:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5370:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5371:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5372:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5373:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5374:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5375:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5376:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5377:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5378:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5379:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5380:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5381:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5382:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5383:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5384:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5385:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5386:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5387:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5388:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5389:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5390:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5391:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5392:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5393:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5394:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5395:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5396:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5397:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5398:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5399:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5400:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5401:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5402:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5403:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5404:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5405:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5406:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5407:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5408:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5409:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5410:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5411:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5412:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5413:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5414:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5415:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5416:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5417:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5418:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5419:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5420:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5421:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5422:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5423:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5424:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5425:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5426:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5427:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5428:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5429:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5430:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5431:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5432:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5433:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5434:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5435:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5436:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5437:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5438:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5439:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5440:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5441:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5442:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5443:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5444:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5445:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5446:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5447:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5448:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5449:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5450:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5451:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5452:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5453:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5454:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5455:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5456:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5457:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5458:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5459:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5460:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5461:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5462:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5463:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5464:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5465:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5466:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5467:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5468:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5469:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5470:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5471:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5472:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5473:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5474:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5475:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5476:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5477:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5478:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5479:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5480:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5481:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5482:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5483:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5484:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5485:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5486:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5487:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5488:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5489:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5490:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5491:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5492:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5493:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5494:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5495:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5496:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5497:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5498:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5499:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5500:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5501:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5502:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5503:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5504:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5505:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5506:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5507:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5508:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5509:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5510:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5511:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5512:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5513:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5514:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5515:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5516:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5517:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5518:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5519:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5520:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5521:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5522:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5523:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5524:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5525:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5526:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5527:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5528:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5529:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5530:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5531:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5532:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5533:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5534:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5535:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5536:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5537:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5538:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5539:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5540:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5541:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5542:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5543:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5544:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5545:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5546:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5547:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5548:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5549:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5550:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5551:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5552:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5553:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5554:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5555:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5556:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5557:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5558:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5559:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5560:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5561:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5562:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5563:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5564:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5565:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5566:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5567:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5568:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5569:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5570:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5571:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5572:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5573:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5574:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5575:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5576:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5577:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5578:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5579:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5580:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5581:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5582:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5583:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5584:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5585:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5586:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5587:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5588:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5589:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5590:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5591:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5592:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5593:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5594:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5595:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[7];
          end
          5596:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5597:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5598:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5599:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[5];
          end
          5600:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5601:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5602:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5603:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5604:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5605:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5606:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5607:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5608:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5609:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5610:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5611:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5612:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5613:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5614:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5615:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5616:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5617:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5618:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5619:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5620:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5621:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5622:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5623:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5624:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5625:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5626:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5627:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5628:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5629:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5630:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5631:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5632:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5633:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5634:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5635:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5636:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5637:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5638:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5639:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5640:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5641:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5642:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5643:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5644:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5645:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5646:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5647:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5648:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5649:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5650:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5651:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5652:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5653:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5654:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5655:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5656:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5657:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5658:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5659:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5660:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5661:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5662:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5663:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5664:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5665:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5666:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5667:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5668:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5669:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5670:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5671:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5672:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5673:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5674:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5675:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5676:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5677:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5678:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5679:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5680:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5681:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5682:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5683:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5684:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5685:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5686:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5687:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5688:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5689:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5690:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5691:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5692:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5693:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5694:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5695:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5696:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5697:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5698:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5699:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5700:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5701:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5702:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5703:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5704:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5705:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5706:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5707:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5708:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5709:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5710:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5711:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5712:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5713:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5714:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5715:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[7];
          end
          5716:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5717:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5718:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5719:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[4];
          end
          5720:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5721:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5722:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5723:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[7];
          end
          5724:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5725:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5726:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5727:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[7];
          end
          5728:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5729:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5730:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5731:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[7];
          end
          5732:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5733:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5734:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5735:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[7];
          end
          5736:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[0];
          end
          5737:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[1];
          end
          5738:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[2];
          end
          5739:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[7];
            cmp[4]<=key_tmp[3];
          end
          5740:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5741:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5742:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5743:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5744:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5745:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5746:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5747:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5748:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5749:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5750:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5751:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5752:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5753:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5754:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5755:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5756:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5757:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5758:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5759:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[7];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5760:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5761:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5762:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5763:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5764:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5765:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5766:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5767:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5768:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5769:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5770:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5771:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5772:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5773:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5774:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5775:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5776:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5777:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5778:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5779:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5780:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5781:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5782:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5783:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5784:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5785:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5786:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5787:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5788:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5789:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5790:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5791:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5792:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5793:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5794:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5795:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5796:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5797:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5798:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5799:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5800:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5801:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5802:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5803:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5804:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5805:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5806:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5807:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5808:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5809:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5810:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5811:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5812:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5813:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5814:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5815:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5816:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5817:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5818:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5819:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5820:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5821:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5822:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5823:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5824:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5825:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5826:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5827:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5828:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5829:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5830:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5831:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5832:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5833:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5834:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5835:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5836:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5837:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5838:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5839:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5840:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5841:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5842:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5843:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          5844:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5845:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5846:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5847:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5848:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5849:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5850:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5851:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5852:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5853:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5854:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5855:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5856:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          5857:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5858:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5859:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5860:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          5861:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          5862:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          5863:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          5864:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          5865:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5866:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5867:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5868:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          5869:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5870:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5871:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5872:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          5873:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5874:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5875:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5876:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          5877:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5878:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5879:
          begin
            cmp[0]<=key_tmp[6];
            cmp[1]<=key_tmp[7];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5880:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5881:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5882:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5883:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          5884:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5885:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5886:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5887:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          5888:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5889:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5890:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5891:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          5892:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5893:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5894:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5895:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          5896:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          5897:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          5898:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          5899:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          5900:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5901:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5902:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5903:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          5904:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5905:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5906:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5907:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          5908:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5909:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5910:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5911:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          5912:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5913:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5914:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5915:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          5916:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          5917:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          5918:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          5919:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          5920:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5921:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5922:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5923:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          5924:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5925:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5926:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5927:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          5928:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5929:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5930:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5931:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          5932:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5933:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5934:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          5935:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          5936:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          5937:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          5938:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          5939:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          5940:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5941:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5942:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5943:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          5944:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5945:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5946:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5947:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          5948:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5949:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5950:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5951:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          5952:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5953:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5954:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5955:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          5956:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          5957:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          5958:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          5959:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          5960:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5961:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5962:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5963:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          5964:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5965:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5966:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5967:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          5968:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5969:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5970:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5971:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          5972:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5973:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5974:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5975:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          5976:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          5977:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          5978:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          5979:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          5980:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          5981:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          5982:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          5983:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          5984:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          5985:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          5986:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          5987:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          5988:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          5989:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          5990:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          5991:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          5992:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          5993:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          5994:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          5995:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          5996:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          5997:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          5998:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          5999:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[0];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6000:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6001:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6002:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6003:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6004:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6005:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6006:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6007:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6008:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6009:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6010:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6011:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6012:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6013:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6014:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6015:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6016:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6017:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6018:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6019:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6020:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6021:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6022:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6023:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6024:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6025:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6026:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6027:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6028:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6029:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6030:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6031:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6032:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6033:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6034:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6035:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6036:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6037:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6038:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6039:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6040:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6041:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6042:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6043:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6044:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6045:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6046:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6047:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6048:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6049:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6050:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6051:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6052:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6053:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6054:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6055:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6056:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6057:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6058:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6059:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6060:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6061:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6062:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6063:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6064:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6065:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6066:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6067:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6068:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6069:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6070:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6071:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6072:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6073:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6074:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6075:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6076:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6077:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6078:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6079:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6080:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6081:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6082:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6083:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6084:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6085:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6086:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6087:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6088:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6089:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6090:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6091:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6092:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6093:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6094:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6095:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6096:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6097:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6098:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6099:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6100:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6101:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6102:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6103:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6104:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6105:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6106:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6107:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6108:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6109:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6110:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6111:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6112:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6113:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6114:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6115:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6116:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6117:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6118:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6119:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[1];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6120:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6121:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6122:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6123:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6124:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6125:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6126:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6127:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6128:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6129:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6130:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6131:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6132:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6133:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6134:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6135:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6136:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6137:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6138:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6139:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6140:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6141:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6142:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6143:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6144:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6145:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6146:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6147:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6148:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6149:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6150:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6151:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6152:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6153:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6154:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6155:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6156:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6157:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6158:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6159:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6160:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6161:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6162:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6163:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6164:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6165:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6166:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6167:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6168:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6169:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6170:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6171:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6172:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6173:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6174:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6175:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6176:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6177:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6178:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6179:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6180:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6181:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6182:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6183:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6184:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6185:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6186:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6187:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6188:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6189:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6190:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6191:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6192:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6193:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6194:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6195:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6196:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6197:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6198:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6199:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6200:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6201:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6202:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6203:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6204:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6205:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6206:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6207:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6208:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6209:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6210:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6211:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6212:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6213:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6214:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6215:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6216:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6217:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6218:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6219:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6220:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6221:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6222:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6223:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6224:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6225:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6226:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6227:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6228:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6229:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6230:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6231:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6232:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6233:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6234:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6235:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6236:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6237:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6238:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6239:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[2];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6240:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6241:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6242:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6243:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6244:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6245:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6246:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6247:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6248:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6249:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6250:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6251:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6252:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6253:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6254:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6255:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6256:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6257:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6258:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6259:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6260:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6261:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6262:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6263:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6264:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6265:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6266:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6267:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6268:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6269:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6270:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6271:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6272:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6273:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6274:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6275:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6276:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6277:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6278:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6279:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6280:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6281:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6282:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6283:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6284:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6285:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6286:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6287:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6288:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6289:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6290:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6291:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6292:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6293:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6294:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6295:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6296:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6297:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6298:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6299:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6300:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6301:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6302:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6303:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6304:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6305:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6306:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6307:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6308:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6309:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6310:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6311:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6312:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6313:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6314:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6315:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6316:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6317:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6318:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6319:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6320:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6321:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6322:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6323:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6324:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6325:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6326:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6327:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6328:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6329:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6330:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6331:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6332:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6333:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6334:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6335:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6336:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6337:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6338:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6339:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6340:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6341:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6342:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6343:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6344:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6345:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6346:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6347:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6348:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6349:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6350:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6351:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6352:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6353:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6354:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6355:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6356:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6357:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6358:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6359:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[3];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6360:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6361:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6362:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6363:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6364:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6365:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6366:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6367:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6368:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6369:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6370:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6371:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6372:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6373:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6374:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6375:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6376:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6377:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6378:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6379:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6380:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6381:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6382:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6383:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6384:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6385:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6386:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6387:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6388:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6389:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6390:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6391:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6392:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6393:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6394:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6395:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6396:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6397:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6398:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6399:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6400:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6401:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6402:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6403:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6404:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6405:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6406:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6407:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6408:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6409:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6410:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6411:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6412:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6413:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6414:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6415:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6416:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6417:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6418:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6419:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6420:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6421:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6422:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6423:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6424:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6425:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6426:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6427:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6428:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6429:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6430:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6431:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6432:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6433:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6434:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6435:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[6];
          end
          6436:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6437:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6438:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6439:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[5];
          end
          6440:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6441:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6442:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6443:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6444:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6445:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6446:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6447:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6448:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6449:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6450:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6451:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6452:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6453:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6454:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6455:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6456:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6457:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6458:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6459:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6460:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6461:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6462:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6463:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6464:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6465:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6466:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6467:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6468:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6469:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6470:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6471:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6472:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6473:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6474:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6475:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6476:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6477:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6478:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6479:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[4];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6480:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6481:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6482:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6483:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6484:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6485:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6486:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6487:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6488:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6489:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6490:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6491:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6492:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6493:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6494:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6495:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6496:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6497:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6498:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6499:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6500:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6501:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6502:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6503:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6504:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6505:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6506:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6507:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6508:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6509:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6510:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6511:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6512:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6513:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6514:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6515:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6516:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6517:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6518:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6519:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6520:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6521:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6522:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6523:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6524:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6525:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6526:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6527:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6528:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6529:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6530:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6531:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6532:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6533:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6534:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6535:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6536:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6537:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6538:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6539:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6540:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6541:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6542:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6543:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6544:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6545:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6546:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6547:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6548:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6549:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6550:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6551:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6552:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6553:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6554:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6555:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[6];
          end
          6556:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6557:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6558:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6559:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[4];
          end
          6560:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6561:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6562:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6563:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[6];
          end
          6564:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6565:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6566:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6567:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[6];
          end
          6568:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6569:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6570:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6571:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[6];
          end
          6572:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6573:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6574:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6575:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[6];
          end
          6576:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[0];
          end
          6577:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[1];
          end
          6578:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[2];
          end
          6579:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[6];
            cmp[4]<=key_tmp[3];
          end
          6580:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6581:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6582:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6583:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6584:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6585:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6586:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6587:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6588:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6589:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6590:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6591:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6592:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6593:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6594:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6595:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6596:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6597:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6598:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6599:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[5];
            cmp[2]<=key_tmp[6];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6600:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6601:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6602:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6603:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6604:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6605:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6606:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6607:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6608:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6609:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6610:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6611:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6612:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6613:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6614:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6615:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6616:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6617:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6618:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6619:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[0];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6620:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6621:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6622:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6623:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6624:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6625:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6626:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6627:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6628:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6629:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6630:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6631:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6632:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6633:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6634:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6635:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6636:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6637:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6638:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6639:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[1];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6640:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6641:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6642:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6643:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6644:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6645:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6646:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6647:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6648:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6649:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6650:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6651:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6652:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6653:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6654:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
          6655:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6656:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6657:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6658:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6659:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[2];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6660:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6661:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6662:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6663:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6664:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6665:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6666:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6667:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6668:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6669:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6670:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6671:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6672:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6673:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6674:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6675:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[5];
          end
          6676:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6677:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6678:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6679:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[3];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[4];
          end
          6680:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6681:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6682:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6683:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[5];
          end
          6684:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6685:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6686:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6687:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[5];
          end
          6688:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6689:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6690:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6691:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[5];
          end
          6692:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6693:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6694:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6695:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[5];
          end
          6696:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[0];
          end
          6697:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[1];
          end
          6698:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[2];
          end
          6699:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[4];
            cmp[3]<=key_tmp[5];
            cmp[4]<=key_tmp[3];
          end
          6700:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[1];
          end
          6701:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[2];
          end
          6702:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[3];
          end
          6703:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[0];
            cmp[4]<=key_tmp[4];
          end
          6704:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[0];
          end
          6705:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[2];
          end
          6706:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[3];
          end
          6707:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[1];
            cmp[4]<=key_tmp[4];
          end
          6708:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[0];
          end
          6709:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[1];
          end
          6710:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[3];
          end
          6711:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[2];
            cmp[4]<=key_tmp[4];
          end
          6712:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[0];
          end
          6713:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[1];
          end
          6714:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[2];
          end
          6715:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[3];
            cmp[4]<=key_tmp[4];
          end
          6716:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[0];
          end
          6717:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[1];
          end
          6718:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[2];
          end
          6719:
          begin
            cmp[0]<=key_tmp[7];
            cmp[1]<=key_tmp[6];
            cmp[2]<=key_tmp[5];
            cmp[3]<=key_tmp[4];
            cmp[4]<=key_tmp[3];
          end
        endcase
      end
  end
endmodule
