//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5z8foqlEA1E40g2nHX1V0rylPB3oocN5exAvx05NtKOHWXqBsAsSWoA2ghdbQGq/
fIDFTCgpSbEJoABZz2KuUWCxd+DJ24vLhulsJNcqO8GOt7tscByTQnh28P7m73Ol
1ELdKAWUZLwRw2h7u2J6S+b7aCS5iU0RzQW/Xdm4yR1WkbbDifOH5Q==
//pragma protect end_key_block
//pragma protect digest_block
lC5wzOADlUEKmlV3ljQc4SbB858=
//pragma protect end_digest_block
//pragma protect data_block
ntjWzmYiwOJlylIOGL+bvCiOiRzTP8evzl6MxHXh4MQtfEmaUqcXlijpjir/aWzp
ht0tB0H40qlXQGFJeRCP0Ga5ctTLfq+ytFxeCC5BfzY9dbCD86FWyO7/OvRSBa4R
bDCi2j/W8iSX/2vuQXy9aI9VKlmoirx0jh/AzN88qIIb3CmjqNAd0zaQMvfjq0Xl
2q03pq2MUraMBATlgk6YGZCA68UL8S0Qfhm2lt8EYcYiTfDYK5sWu46YWQ3dflMY
v8FPunu/Rqubgi5BcjkV1MEuQjnvTM8qOIwV4iDhZZnC2z5ZxqKm/xSix+Z2VZNq
HZX1fnmFvdXMp1RfT//Y5w==
//pragma protect end_data_block
//pragma protect digest_block
JraMzpUXa4kL9S9NujWsAUZuIHc=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KAhRQ2/mS9P7tAnwGkCxLiKZH7vAHsDiaSGm1fi7FQ8dgdPSNa4Cz/BfnovfLBZ2
OnhYirecUAgOAYGXD1M5imcN1mzYY7FS5MWN6q61M08wpjYlPVg4QE/cwZRJcgit
m3Jmh7oj/WJgnF0IFsxDrPyPyfosualwFieC9VXwF+dhikRdtzqH0g==
//pragma protect end_key_block
//pragma protect digest_block
W0tW8auYb8aSVlM5FalFYQeV64I=
//pragma protect end_digest_block
//pragma protect data_block
7J4hF/j4/GGLX3fcpRqUXyYQvmnYIxVLjZ66c6F4Wgpvv4GQX0fAMLbZihrqTINX
LFG0qxTp6LlcfsDyzGijgUjW0CWzc7VCBNn2hQddHEljALr+fz8qCZwjP0sH+0cT
yTX9ZWaKBfcVyrh9Ygm1eDrJqUbUrPgzJhtGEufY6a8/6Bx4yQNr4QU6Je2aeiiP
DlThnRHCX2jvInGV8NKtdXEo3roXYWkGsLASmPtlQYz179GKqRi2mDC9cCLBfzkx
IpImPbsbhgo5ONNAgEamQ4oW/0EovIWTiovP29qndTH581JFbOGWr0KDKOxRvjE4
sjabpvPcksIrSfWrJvzmPQ==
//pragma protect end_data_block
//pragma protect digest_block
GJjIM2ycpTe7ojj06pJBck1bdBg=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
mEFrIpa4sah53I0EcEaHZJmIlzi9WVMXajnJSAKRSPpbSyd+Wq87FjJfOnp4WHH7
W2Hv9vAsAiiMPr7edB5EYRt2YVKhpQpqKF6gSSbJHHsZ5iC65NxavNI3X/SW1MHj
khRiH1XVjfGFMgVhcKTvdR7Ju2g8ltRYuJAB29ucDyQ9+hZ2qvJ+Xw==
//pragma protect end_key_block
//pragma protect digest_block
j3Hh+2F4ieYSBG/JMufGZ65DvZU=
//pragma protect end_digest_block
//pragma protect data_block
ENac99ABEzIp+ALcX5QbZvPY9gVPneTUy/z7GAb0NnKNKyP6pYoddNLIMMjLQKhU
yWLCLw/09lVWeiRF1iJewHyEmWpOjSq7lfH1zthGLRRFOIavFJkXzQY8b20KzE9G
7XPgpk3y+PQYDaXWiiUjVTjjzbQHGGdrej1Ps8aOmjrKZ4Srd6Wkmm2OPssPdXH3
ZJMw9nNRCSKdFNDq4TTnffO+V3bK3VgNIWOUWddp+4Mxszf+gvqdxXrJeymb+j8Q
hWsnjL8LMIitzSCtdzX00Kdx1EKklsBD+aNh7JkFOYyHx+TRrtChRS85rD/IcUhw
Uv3LQIkY0N4EbHu/kzwUyMediDavmXEaNlSVb6GQuDHx7PzCRBVarqYcKwpMjpFO
ux5AtaHBXaIDeuf+Ok28xSII6UTCKNaT5dBoUXfwxZDdLgaDIxwL3FhTz/0Poc4U
FLNq2uEP6Cg94B1wQxN4tjH+PP8cV8bmP6Ucn16j0zTZjg+Fm0WuG6kOzTM2s8/j
w7LbRu+uR8lvHuS+8WZlGNbJ1Af8C1oT6Vm2enoGHCMjvfDZwVYDTMserA7IDHzg
DMtdItSe2fRt9M70At36F5y2k9A6gesGvNeuwmC0yFgc+UHYpE7UlxppxGv0KSVz
8/PwhwUaC2OQTEMraOyan73C6xT7c8rnZ6ZRs6RhqFA0T8trBGW7cN8LOLupPWcr
H6VEJEM80gvkrajaTkASpo2n9NdHvBPWzKFn0oOCPVgCLn4GgtzqO9lFycR8jsFw
x6flXFApfOmPZv9Tut8IxPhe6lUs9zr1HULqpTJebCVRLQbY0EUOeNQPshv7McS8
rQd8WuhsJDtvZ6adH0fQoruQjYoOzjC/xaAcjCH1YZKlxmS/cxCCUVS4cJfL6zWi
Jg9csrESrRDRWnWOQveN6sYgVCR5gCHJHUmQ4PQoNjunoVg9BqsAEmgMWd1cFSBU
tGbaCCBO7/VqBRFtVeOLrItNQFrii17FbYWofi9bRR0IyTcDqt0bFFaxis15MJVK
UwLzEGzu+7gsYusz3P03/Fxutb/w42vf2CE+i0tcUpOO5nACtiPIqRT1RaRaijln
54BtgyOhnTYZie2x46dJsFVj98QTuFCo5/Ral4sDDWkf1qyecvr62Mq8VTWRap+o
ANlCCDbeSCRBGTPy9r6Ou/+kHQ/Bnnvm2JLSzXwDfpHXabWDMmJRqln6yRBasL6m
ggXCXOY/8ruzbkcvyns7tY3Hwpj5t/aeUsUBACGDsLad2McFXKywblStOaQoF00O
Tg+ve8vNqGONolLDHvS/szMh/HkdexCOhcReb78o+9GeCkx4VyZkP1mSyAC2e+eI
5tkedQDglkFmrv9qHTmywkzUwRkn7yCGeoJOxT23I5ewP7eUPYXgicyf0PEbfgzH
Sywrg6jBLc1px8lAJfNkxft/WJ9QAqDXW5/7tzgfEIpAOKknrMWoz0wCzn1rfDZ2
oaYGuzWI8ua6e6gh7rH1WRXPnsgDRdIg0H/Hb2CF1JxvC/Mi9f2Rs0VhfCZ9zhD9
oDSihZCQwfKVILW4H6Cr9I+PlAhG2RhxDjBYjsCi/WqoaSSOv71nlWlFbzrKKH3i
XWeTa+S1Uc+M/LiULVBsO3dBUW+Utx4GW8ggeZUwJrQMDosd8snLeNiJxKubbLau
ArpFwbp/C3vVahGjtecq4HkDnXW7rGs0UCrdA9wsDSZbz+4q4Xm1d3s3GSrXLGMc
QhCjCIlRn886ijt57gkaMfTuU5IwSo5QuRClLXJX33LQ3lPbePUQtdyterw2nLu9
L4UF4kxz8ADQ2jidhNpQXfx+okQ4dx4P9J4mH+5CYV2DTJpXr6ssGSVrH/V6DxT6
2sdgx8kmVD7zunnt2hwi9t96lE6yzvWpg1CE1NK57Ur1yWoXx+vxWu5rPEcC/ZiV
F27mbHQsMHdaZ47hzpUex3Mdo1UWQVmiDNxTWIIYTfnOFiO/SHJ5QVv/pf+EGyvj
H6ei2wA9nqZj5CAW7Pq5Q7qWnGady2/OTBswRe1LD9KkbJhRTuk7SgufYvIDUCJI
dqbh3/0Wr+3gkWRXn76LNeMPsg+75uvThMKyOGIcAHKsITR9hP5qj3X92qFHJd0b
oxsoIRYCoB5lVCL3uzZanrvXIej3erq6Cl05Mym4LY1ttYTtaM+MBdRyM+FgnesZ
9LwPIw6KhhAq+Zjlxr/6yai65YfZbeor+9gEwOPUwYOU94xj4kg8jjyjlb6AMunH
UMNAusshiPW//DZeW5RT/L7Yr+jmKIeaz3IVAaG1+xGsYCdDn0Eoko93+4heM9ts
bg9LKHQlLthfAOazyoeAVIqTB2aRYG/6riVtENVAsRntg0n6wOencCAvOAyQdfa4
v9Bbf0PhqQZLIpMWssqSkQfSgPAI8AuVTaOpon5gk6bwzms5a2ptq31qXPFmhnlE
hYM2hz2CsaXtZybhiy0WzDsFsD6AFmnJSMrpKSTMnm+FtO7GYHRM4YQSWZJboM4u
5A25okXV/BLUcQF3NHbArHevLIG114us+rwKDha+E9XkfOJKxJ1ONHJAgHrcE2NG
S0REGZd6BS6isIvrDGnngxukb9bQrDb3C6Gc2C5VxwM/yIyaGkq9/o4Qk3+1j3E1
nh+26mVc2j1cSl/8sQOqJ8CzIwsnhLH1xt2W7j8g+rXJ0J9te/It7FIPhZzFU93r
wxHc91N/9SRGbxU2UpnYpzOy0WKk3nyZX0h+XuX0rjKh/0qOK6giNbanekXa6qOP
bOnFjD0ulhSujAKTp6dSvf+6eYj+6fMawxFKZoysHYpOzBdpT+ORkqLEZc89oWQf
juK6WpnUx5B6uI5TOOXOnI18e2Al7654j4Ns49B022EKc+EkZMti3eURQWihbpVg
g65umwBMTX2ERZQ2wAmA3QflWLMLriKU9KAwH4HPeXz2Dc6oib/QYSDUA0oAqQLJ
EY2pT1RK6f8ZXsNoqW5BDYgSCyvjsQaugMHt8++tRHzRu9ZZLRqc7nttlmo8RUEe
BRSeMaPQGeKzm7M7mrrsey8JDIhSeWUIv/Yim4gvd9oz1QExhslFxbeJGJfAt0Gl
d4/YmUDEuSmDRBC1rUf/1/VNzIC3nQ2HN4qcODCt/Znk2tN8MjU36fC84ABNXe92
bY6jXStj0vxHOoGtFZsJXR42StYcNVllcZ/tJpOUO8ltdWzoPomWPRVYI67cAigk
QCEAZR0EncvSj7NOsR4Oafdgf2hDvNBEPT4tM47pBioall2IOa6bgnWRP9GIuNTX
I0v+thMFvP4bJ8H/9sGfJhT18G+aJzCyJfCplxpMtgsLaiRbCnJK28aykAoDYgaP
7VA9g8eUUS+aWl7wLVJs+Fzg2IgHuRce+iCSUw48MZw8+OQRSL24JrVq9cMiyeg2
Z3MljIEaJAqmqvgl5VfEe10fTR7Y0gQqDB6OvClLK7Pi8E1XolBlkxeS3XOwgPd6
+OnQHFAorjS65zKjEirUR2EOKKqDuj+Q8LfAP7E4Vh4cNCOBzZyZgugAeNIgdYR4
XlbnspgqGsizZnZYgeGOywwhgukhf6kn9anaV5CCOtwyNS3ktYSSLKRwfN42qj93
w2O9waZNK/HW8qC+mN3B1xH5ovA+iohMCY2I+Dq5UTJsvny7Ajj5Ev4NPl46khWt
2hT5BI2i6q7y5IKdAwf4nVWc41oozdMjlE36ETMC60DDlnDdWcSBhEarPl0xj0LD
oAZsYtawcuth3HPNl/QfW5e5CGjgJ8+tbZMDukZsiOQL07t4XNFLtfzdHN1XVImT
HXGGVaxWduqBChc2qAhxA0Tg2+6mJ7JLUq1BStXPwBue389Bkv2rPcRIDwHL6Z2S
MOzBqsQ9onl7F5u81Z0UxxU0BbXrj8Ep8c1/dDUwSfuci79/bszBe9ywMIDIPPEB
7mENg7nzUoXbhQBFrYk+O8ZkKZ7qtjdQQdDQYjOm8KGuSasjmylcO78ApsFi7Us8
2/YHvN0XDZbJgoAfy1Hyw1OpEzS7izsLKZzaFJq7m9LI/Lt1l96DCamhZVwOQ9+z
RCWJ2oKBH2C3JqZsSfh9hEeoxlwQcKJBQRHLCbt/LElL7GOs5G2VvNVJ0/jnLG5S
Qx6YXOOMcAhqEmleZgcee9UKswaJ+hPVLR2t9sK3iiaBeQ1vSIPBgiUKLRIxcvQv
oIww5BLBCzxhJOy8TByV0WZ1C0aYrdopLIz4ri0Zfr/jM97kbdjBHwBCfDmbqJhr
aZ2ZEzmhfibypLJuzsX9W6mlDACYpeeQ6dfkyJKrNIusoRCcecbVZBuxSIyohr9V
sIFQ5ZSM5OWtXGHc72TxOVX7zX4LsKjkCjet3tRCmIQQvBH91pmETEfS4QnEzgdx
o9wJGGSjj9QEgKGqaH9MtShuRGj8PaAZbYcwfuUJzefGvHAJ3FHfCPsyCEVyInr7
tB9hQNHpCopc+91Vy9wdHsB61PwzyWMWD7wduvs6DMW62nEMJG10TEGoJNfpQaja
7spxYiK2rfdWnb6gZDf/aMR7cVTlc6OWPPtkxkPpS9b8uOv+IieokUSt0wDw+UaL
SuafufvhU3oARUwGLsZcuN/qqsso4I01c562v/ZskslvBw0V76szYnH0qkoQ4n0B
WRBR4Zp3BrbHV1tVCm6J/Ikn1WBpsK+E7AeX5+UEDbw4duWeIov7gYi+DQXmEqhg
quws1TAaY8Sh/koU2R5gwpLJuaDfHExYtqFUCajkCOl0VU1VHvhXYV9ZDMO8gE5v
cfk3e8KaUh6CgtXTSGGiJUvIEq0YtYKWO8P+ypjc4U6qCzetnVXNzQv4+6LRSnyI
9oq02JCfdgPqvdijZpUvUsSzu7HAMGp5nyJCSdejEOIEFHFud4f+uH4AF7zvP15w
zCC71jY0DeUIFjY9itRD/FbDaqdI4qFBiyjQcKHgi7+q4l/Zhs3bG/yAH84rT0AQ
uBPKuiRZWhe4M+QogvFHByYnUImAucu7syjYfDxOXAoFnqY3OCGR7FhmqdrzEaez
Hu1K/6lstYZkV0at15Wn6XwbFbdNTL9ZnqJ8wovuKLzqFStqQw/hbHQOdxeMiQmb
JlBtCcoRx47Dru9pdWaNVWJM7MRQygIDXhWOswKz8pTbWsvaEDhYRRMoQORumpkZ
bv4Eid8OdexCots/ix8+zhG0odD+ArMZaYEeAhcM6OI6lLwHPlQ/ro5c6GXb7gyL
SF0G6jXLObOmCrY7DEhCbkwcbx4B95FpTmRl/pFwxlgE6NNZUHnkgdi7yBv5DzqQ
CU4e/dAMNC29QPJAxr2djTEUue3izOyBXlk568Ygle6zPyu+0RJu4DrudYxnV9K9
J2FKrXbxwNmfuLDTZ8iTQThwkYEnazouPmpyo7kXpIQo423RfGKzLF+2Cnr8/Iso
m+fBtWNMtg2hUm8eSNwI1Ryk0fPKOrxsn0L+I2LDWYbbMlk/O4CyPwGSTBpsIe5J
gylUkvCdoLvNajfydj/ZiOmmYXfgOUgAMAuX+z9zT8IKMTVR/tqQkMzG+yyt5ort
2ZdKbjglykSI87XQSKMTuu437HIUMZxGHvukmZdNx8Rgd0UcbOMMgRJRVH6ic8xe
3F13Ef10VWqKVN4r4Cpb+yNHXv1N/GVu2j67MFB5s/BYGfsBUqQDe5rGiuTk47Lx
WbN4IiZGTsknP+4WGXeUv95uQnAGvJONTOBx80vfM/J2Cu7s3vowpJ89f9m0H/gW
ACnmKECeRXE6ttdJ6THRghSIexrrODhATvB7TsPfewjgA2S5DKu8pN/5tbQUo004
Ll8tXo4XBjp7juLHATigCT24UI/oz+f4tDKhkhZpMGxbgbUxjdWurt+kW8U63eOU
orr4IQJJ4op4/kvLHFoo0BwvBYlmfJYMru4mFlW4InRlW/DIaIvxxfa49mo4KdEO
UJ96YAcfTw6BERHKt28NWzuVH6pvM+qkRgSPph45hA4gg8P8AKqbxTLguU4zKfIU
ejAgtXgFJYH/8AzJ/lFcDIlh4oMtRl/Llve5qWRXfUk6g5nTIU6dXZRIJ6H9Eg25
LNO7v6PByuYH9qI5PODbTxii4nwXJrejvAEB8dvgCiUxq/j2Vz8P+G4o8vdWVqVC
TfJCctQM45SXYwgspHJiuGbafheeMIwEYWPetd4sncvQxv/V27rir5MlKqr08fxj
fqqdFl5TmXubSSwnWREsMl8VCz0/KMbQVjNCSzDzEke0GlQ38kli6nkk9j/XPjW9
eGOixpPdmz2cZFXI4uRRrdIK/C1RyF1iHe4AMKXo8PqQNNJbpggQqxut9HvrrtCm
/qW3IzLGOJD0CefMNIFDZ49tPLHnZhxpV+dWfCpVA31224he6ARmiMIguqOCJ/il
WPnjPUgd1/NDAI4q/21DFMftw/HjeUztwZqzA5HxRiR6iZCq4brem8noJ53DUjGe
JXiILtJbtBiQWtFoGckTyXYzoo1zDVi3u2ZZUi8KsLMZGGnsyG3Z1PtTsPG8ynpC
fZ2Z1SkI3g9NdZajZHU9M4tedEvl+vmNEtdtdJ7lS9+u0rIDdp2ZV4no4TjReEdd
i5y6UczfeShJr/YEqN2EimTvQWfvOJnewVMJ+K8gOvZES1dqpPbX2//Lk9HgNYNJ
TBGe2/vimTv+7dxUkDNumXXnYMSbpAKf3dmPtmViN48fp0j7LQ1ESLoFGm3v38Iy
iVQTLLXCFGK00WRHUP5ixv80VKzOUbeTzhO81Qvzua/wf2gk4ZjB3jRnRHDav3QA
90knNerpK2AquERWUohh97B+cD0Q26YpxY2mhEdmHhhx8vQ8b7Bsodvcz7cadHa8
n1GPC4SgpT9uka1NnDXEcPBjnhGC3zDZmmK6mt6Tuh38MK8nAPssrhmayS2OztiW
+Ab7YIEDe78UhfP0+vpN84vUS81xlfBIqEyRLBDk9SB+g0h5zPVwIRm2Yes8WsmY
sIGnO/xYjFgzfAIQpM0T7eEwkj6VDq7B+TFSWWG7ZEVjETO30TpVknomHAWO0krK
L8PzluYXW8lYdiwxCa8/6XxF9ZbgmLwVyzkfH25U+q+00KOLL/AYt5xWLPrTLmso
8BPL6VMYD4ywmD7w/iPntWvEu9Pp10MDCE16/Gu8n114arviz3C9eIWi0uZuW54S
EhkvmKzrHQdnXjabUzXDWNT7BBQBVP3KBXLFX9JE2soz7d2dIIbUcjJXi+bIcgcC
gMWi4DEwL/whHTIUNPjkqUMK5UYeyaFN2TywW7nyFN1shVQ9O746eEKY4+jnttf2
hdr1Lciqx4ImhdWgaJotk4G3x0lhUWcBoK/wwkN0pXdcU3tT/sx8GPYxgqvtHccl
afoaJQpp+ur/wumTJd1zxTGPZN5l+/7/VNltpxf8S+sIU1LvixRkgGwZoU50LQbb
YUcyMgAs1eqQ+S1JB8xvL0SuLgfoGAxqSmn/gtYlHwCKrvs0ZzmwMY6bdXgz3E/g
j3Z1Ma1NBL+kHnH7svStkmdIRLa7ZJQbt6ykBdOIsebiMmvxGeMVJShlgk9E0tIH
yqWNkgC75VWsMZEwuZQuwEDwZ5/YNLL+ABZk74a4EZT+rE4bZwLjlxeAVGEi7bGb
clKauT9QkEQ5XsemrJbMbU783MNwEWjwc/UYOzQJzL92c00cS1jEPltTiD61Nn44
grUE7WCmAXpHDjNdkapq6Bu3gqZzX+t6ealteQ0B5pBgKDobmsf7rRWvA9vRz0nD
elpCtmSZt/s5sgRQBFpKdrcE6GITLfKnoaFlbjKqc/rxIjp1ZHqGt7CxNXX2Nyy7
RyL0kD5si/+QV7Wu8LLTK1Xr7fLFg201pN1LqctIMNClXOz2S35G4lE6YHPqGFTV
kShMlDppKjXE8FYSnzArEidPrVO5jZCRkXullXw6924JqDiSRkZtPH/cpkdRERWR
QVptFCKPB9Irflp5kJHXBHBKzuMLre3Q3cD9fcmUNS98BSpk5+s9OSdJXnu/VJMU
zgOpWyJxNaVAwya6fy3GYf+oqXN6Zwob0MZ6fsFVEnB9WyC9g3TMJHO23XhDdLTc
gze/pofaJugAZ9H3TFVZT7Ejwf4AoDBYiLlYCLrQkI8Q7GNQtOPE4f/4k/rpYmgQ
87vSPkVdj0gjzbO63Wu97bYW1MxXURIQx7ILaX5GPqfY+k8MTa2XlcgXvWEY/M9I
uuvpjexrPz4pkFu9xr4KPKB9joG5zqxahXlBjZWuK20s3CxgpYlaEQmU6zkqSzZy
37HLrm2H5UBX9+85fK4q7YtbIkxnuruT3xIzOyIPFmmBGBrjNlLCg1ai1vg0Gf+4
yxIhh7oXbXKdw3zvWif1MVYnS+lEpkmVxeI8NCcgq5XM0ejX068An7V5M9q2SJ2L
IGSf55ETq16pQMqUYe0Alw7i1xFPNL9SCVRleJbie5XI0Wdgoeh8Q4LFxyYF3icx
TDQpPzkalI+ZNF7MHa+fIdwMgdan7MUIrimIP/xWPGVtCP1QlfwX8MJvzdqxyj46
2a0D/BHwJmDkJKMBLril3kzE/ML4vpZCeRXo6to7kFF8YHeXUuDsUw1lXC+tKCii
z2NIrWTYp/l8Dh7FqCXHDIrNikxnlMzo+VMOskiuoS5TNmzcP7s7W7gukbgZJzbC
szVKYC6RL4Sg/z2JejFw6z7C4z0cq+zjuOuhgO9JaTKw8QOQsBWNCsVo2vq1lq2W
zhLvsvOey/jymetMEg14fygFYUPiLmLINLzle0DepZ9Bly+zYhYQk0wQf1eN0g93
hUXefG1ckyAgSFslG0dpmE2saEmAdAQIwHhMPEE7ZQ/9jtV7+lDJaeVtnX5q9L3H
3j2Yh94tG8pk6hjZLB40EBuX7JwnAIDZbpzww28Ki48+aYJXxC4Y5ZaWSTfWM7gQ
FUo+XxAokDTgbLPb0GaoWocbWJwWWvGMHKkVFagOgJmKf6u5CNIR6/dlmQMX+9zz
yF3zF+oRrNJ3Y1ciOwnDWDnhiM898t2bMIc9rbZNc2FB1uuMYCHqoGcFYASJuX2Y
l6ZXytYWsgik/UQbM2A3tKqqsWoTOgN9fIr9J/K+zAKjQVLLUZc0DEQR55vYRN35
yUG4JChHPve2jiJ00rsQOKx8oNCxxuglowANfRAbM7vzZByKwP8vyS5OMw7zsLsJ
UYZOE13VP7hj8en8hDyXvDas5RW8K7PUxULqvM0+acWLqD8zVZ59U366E2N1ECAN
DgNpIwgXIU0b7Lq2r4UTK43uzNRO1y4RzbOBV/y/HByLMVUXOBqJP77kvKnR236l
TPf6ivkxjmCEN6wP/IDN/QgYZCKhg/7G0WbqgLLVZq89bjGsjCrbFTpz86wvF1PP
c+YkBOGTokkDkf3G5QashcC6o0PxVMwyuUefNromW7lpV2pX4ka78N82vknJMTKW
WtnA74I5k8Y/KJbRrH/tKPtDERd6mH+QXdVPuH0BDb2YqtNgQ60KJPefHW6u8Kbz
dcXvOHJYh6Jv7ICeX4yVpM0hVxEUNqK++TphcO9KrVq9dAkmwtgEL+Ayq5F3NBcf
qxWqJKz3NefiKm2pTW/T08xxqQXqsN3vo1OX+1Dpy6T3hvZQ7vEvj6tQnisSVd6H
yH/svHDv/ywOJtHOcOmk3GpGpUCPop2W7pycvSa0lPDizxCTijBVmPwPHXL8+Zti
5XVuZbLcAfgB1gBe3/cyHmAoyu8dyCLobJSnhjcw6ZumWB8PPwI2St9k7YoBKgKA
ErzVQeq+xOAp7bqnRMlbxr98xf/iAtDJs4WYMBWSrOXu8JLSw6UaR561PFNgheNf
1tA7ThWKgS96auK+jJCKxvIBjrHOc2G6klVQ3NmuyigAnIT75gaaQUt7qGqzizZL
vRmqnfby6AQF/bu+D39oxLn+2Y1vh5REJdY1JN6LkjC6qYXp3I+3pBk5kiGaNBJH
cFLaBMFGgbBWDLglnKSJdgP+1ivcFFAAeiBFO16PkGJqDtro2cQ0j2Ema++1qHuq
4Pbbwf+DMecw5gmR3Ddnj/wLVwO9bv2xG+7I5aPKxUmN1xgXTp5Prj8p4IUpGzm/
TlgRGI68wHVp0t0+it5v+0eMXQ3CW7V+jhLyrb4IqIki/7nIpWDshiDVsfGiD0Rp
dNnsIpKXFbVLtAzLDlSvrFn3bieCruOQMtwuRm7Rw1p0hj4zbns263YUWlfnNg5r
oGnMLkjwMD5W/xHNB6BlKzwkFbC8CJtKB+vfSISUJkno3wcQuhCA9YeMM4hakViQ
GlJrd5jyWfSB8ALsd69WDQpwlYjeQ0e7+NfHub50jlwXG8dFWpT42l1hjPk/y66T
3Tba1Vcu9owfDvqDS3NQ6DQ15TJhbKDX9kziTFpyecGEysrypu0dXSsRzKzW5Z0E
dMXsjnvyURK8/usPTJeGf9aXpz5cBR8QjNL4adzSBTuXhRZNpFh4CzGYaj8wwZZn
jz+FnT260P2aCnZUJjAxgUl+oFWQiPZysIu826hjllLq8AMpjzWxGUFTGL9mWw75
uYt9lQB9qcBwufwbwft0456kA3BxwnYE7syNrIuSJsoiELaKiF25hnoTx2pq/6dZ
zK6lAknkukR2q+dFD3u/eMaT95QEcWLY2SwE1sUc3mJW8eYOOJmTRJJ++/cL2BBN
aovb6Lwzd37k9rrYkGVI35XVfyZgm+vGEBeuIeis0N+10FIB6uSCGl9i+zKrGAdp
N3RSUGPAoWAHAIc73tI9YlfeLmsZXavj8mvibJupTzC7E2l3aRTdsaYFMHRncMon
xHlRD2Q/qnxkIujj5DOWQjuPKFKK5tYV2Nf4Q4WIsOF6jD5wiK3dpGm2tgnvudce
F7MldDpVGNE7g2/SVDWzFjV94XiKxrxcHPKP1Bxksr9bDBVl/PRBpfWoXIq8LVZj
zoxbMX3VHyKh6t2rFcWeROrwTOxv2I63CmKt2awnxGnFBZYF87ldPKDPkwVMaBFY
jPFAXR4psWnbRjygfgqCEBmkwupUCxJQ1eRYa7/cANBIea1/jJHaqd9l/c0hVaWr
kYHM/k+QQHj3Z7pGQZiuqYu2lj9fY0uy0VZmVUUNnEcGWxpvNwInbxrwnW5L3XBd
Z9fkGMbey5XSLZm1HUufCQEArG5+t02sAR+ur+Omn4sdGz4NTft8uu3c+8/YLRmp
vPNMkR1xsb8Nd4izDBbvaD4sb5VYjHIwb5ZYXp63prZzlsKZiCShQkKKttrQdSbn
NipgQ+9J900on2Etq9zhEQw/F2U8hksfjQ3e+QXnuk7s9i74qI2PEvBvqZcGhEsE
LK54AARLaVNIrQ01jQx7qc0HerbsvLo3R+SkYQOgAvsG5GgoF+vpewnHgpPJFuMn
srqtTv0ieA2dtX2kOwEcstY2BVh/+N7b1ocIefn3bzaF0Nino7gkx7vORT7MfmOd
hYIzjhEG+2ajaGCIdQYcIU3pVPzVkGQL7svaTRwwzjrNpGy6AdPjliIiMJzIab3N
p6hThJaD0i3xLOQ53kxQgBIpCokKjYVFBv/LxQYZVFA30A/cSlWT4zlZVHKmQhRH
BjtlIl+WsA8leFOrWmC/1xGODYBBOoM8Dmzvb4f9NXG+FO/8JGRGOGhC68v66IiU
KR/o0AKQsQkbk1PE7CACXBngtEZJqT1LEJR3HwFtnbYo6D3cmx7GoSTRHlPwUCU9
k9H2fK0SXU1BSZBdtZk84Y8S6CbcD1z7jwNj+TLWriTLNRtWPU++Y8D3U9A1Ax8k
76B7466vbsZcA0U+pvOg9gRyPEGHWZRFSNktku5s5Uu5fQj+XHplBibKQmE4zz9z
frfRbQTmip0oPTjcDQr4xqct8R3T+XpxfZ5wlDW9tIbU2K+F59RvB6A7mQIX+ibS
PhtyvajINaViSaSwB7VbPalPjRpebdtn0SoLbAOwEyGMZ7J8EPoxvU8xssDB72gR
7shfpVYeibwAGBsAPKsZIlo/vOriDY2KEMwWxbJDDh031P71H9RZCZoduytTHiec
PwHvx7vbCrV6ciHIIWWtvrkWTI1PMltD76+Hg8SMWudJ3MgWwc/msvIiUcphx2Od
H93ZYtiCczIhz9Z9cgP9UrlZOUfMLCRZ3QBmqvrI6MedI5D/XfasvPvEYlpIuJXt
v7NzTnyLppyMPB0NPQ/hF7e/hBQRelx9VOlAt4eLMRpw4Xf2a4/Tojw97lSiCcEl
Eml9D4FBKvgc8fhtmsrtGz0saUH29F9vp7yxJZtIg+ukHHIM8DEn0trMxv7Q4pRg
Q2bNciK8dVEgDKY2kw8fjzN6XZT90pp+dMY3FhX5ePgiAvnKmpWHFYQ60xsHiVJK
G85w2JY8rd/MFwLtW5/rxZo5bwWGKUd6HUwpx5ris7yRKIwBUJgEFCiaDBGX1JR+
eLVyTMNtuKzGYoIBXwsVcQTNeKOrqE0P1iuQpxkjEWK6EEB/iPvi+4K14vTeBPM2
rbzZPC6BjCxFAqA52+PXGaeS0l+zBPbsWiMBDnEOGYgxRnflwrbaesOvJhhHmqZM
UZ5QfnG8bF5rX284sk5/oiE+TkiEpBJ5RoDN0ojptLR7DN/ZkE0Ed0/byXGnuw8+
F6XAx3NelCSLWK6FROrGCasCSXPGrp2Suqi/2qIRzVqyFrbpzeu0rVGRk0SLAm2W
LITKwIqWf5rrSvAz6UR1ca9ogTibHmX0QRdKSj1NpS6R5StXXBG0NklZLvWSmIxM
/rZjTqMFsqzI1mgYIIRIDsFus04kMhQJYSwprtbOZ+rfF/K9ka/p1YWtdy0MK7EV
/KjFLR+/9/2OvAAHree4QyDlvUMmI0kKhvllyeDYD9ViAnFM+xemZR3XcCKVt8SA
SONK3WOutTaHdov/Fi1CAzvRo/IZi+/oGQeVwl58i3dabTClFDCsRj0UDGNnVMV1
1/GujKhM5kV1iOHB4Gs7mOcTvahNnjG0Pv0c/nNmBuDDyISErxv8rDSY4VwTNcMn
hGBxAW/U9RWUKlaOqGDYpZyWozzJ2+ij/41YKkOFT1h08Gg7QUMKUv2hBA0zzB35
kre3/e0naZVyMWEZBKn+ur6VJUr6toLCF/Rpy++2Zk6ZYjcjU0S7v0j7W1O3PB/K
FODZtNlckBIdrBVNPXngsOWK1eHK36tVYNKehijQvJudAXHm8FiHpIQA/z2mEDhE
UyhCsBqXF9ImtvonMtGxdAeH/0xcuScQ1+l5lfrctUKsB0oleRIzD09xv4WkE8WA
gOb4x/wqaRPN1h4hEne8tgkMCzoF6C5OLIeXJa8I4opHKThwqq2tCYGBtDR1zgjt
tVJzv3cUNDoO38aFwEJwumq8neyCxcYGO4CSti8Q+IPCVI5KVBJoesxr6lcFY7yk
1hQtT9ffoLM6bSOV9uzNO9ikgNj9wbJW06xIzVZRyafXaK2ljzTvPuowfr2Yvwlx
o0uUJhoOfpHpSK3dtSqme+bqJUQsiWTqGoS+NTn8yPnKEDVWgShlthXHfaYBv6p2
rk9J5lw+QjFB3/gET0cfQv8XsTxbcb/v7+DeyyZsa+nk6FZzE7q4DHcnGxuXJ+g3
6YB7seq7TsTV7isDdAHY071RfoCbGytM1a/VibKJnAMx6DK3Uekqvhp9nHU6vBAO
i8uMQ5v9H1JkSo+a1iFV2d6llxwBvhn0jBO+PaQQTGLFqot/Zj57cFO2uEeKPPhC
hkf2Tdxrs13ivWRgJA9aCkQRx/i+PeVA/KKB7bQcVi/xdwLndwkhtCVT9RlCOKBI
AREQVVWu3PE3UqOQPsYHPCVsqQIV8XHd8OXNklXWkcb8rOkTqkiVI0JiXCgD8hFc
oxQTygmYrxtEdLolfbJUnOF46/4A4HWqRRz1mghdQYRSwvj5FcZM8UEX+Ip3s6rE
BaZbowH7deyj1f5WotwS+e2hewjoyGb+4zDn1ijqObaPjUL/0MMlCcKeeRUeYdNR
Px8v5nX32g9GvkaKmV+EJeYi3d0r2R4D33duvE2uLsiPWtcReYClvms4QzjZo0bx
n7JGok+rR4Z7bGbkoZk/GJJXf56agnu1nx9d7U9VZV4LLZFd4hZSnULeo97HA6Xo
IzgsDCnCMmCx+TIETGJthvFFyedLUpqX7IinikUdNaJuz+muesgdw3dcS0Mn70X0
jx6KzIXRJKBKEtbLUB5kVd2T2oxzFALhq8TlwyMwGGz71EHpKN6G9d8uepJzGrLq
5PGkt/4Kddf9OaoHOdbtMe9PgvGO+QYK+e28RmWnSLVyPHC7SP0WBCvrIA842EL+
9asbQ5aZKJK6JfrA+s8bBRQAH/0RwHKyHMnz69IFKv9duwxPERXk5MStSHdxOOw6
IuSTSK+rVS9PqQLWZq+xrqGk0bMXXNHOfRep3XZxvGD82gdLMRWin92lUSUoDv3E
FgZYe9MNSPmC0hMG0kUf8nAHrtH3SMLo94RG5ZCCws/QptCrlT3Zr6NIDPts2hqU
wyXNl7zhYx8JZgQNmH63aTk5PIlAt4famWV6CM+4hncmmy+R3WOx6KS/REi6CXTt
MmsBBmyGdoDswRz9K3TuctN91ae0iJETktlx8q0lIy9TTrqps/U6ybhaLnPX5q80
mEyOTkWdFv02K86PV0e3W9n3uro5KGKsK99J00/RdbmODbyy6z1HZZEHYprT4hn3
UoGv3+ANoe0wdyBc19vMK/X5tknQpnsV3wDcqOQs8llVLQvNJKXllYGwFlvdGfKH
ZfqUnbBcjZHcrRvJIftr1K0jRoyRys1mB8Mf7vXMPnhiTnXLejE6ttItrY8x0yG/
3tPHeGZbfjHMi1x2q6I4puBoP3TodPpRLvg1Iw8PPLeGoG1BzxYGfyyCMsJJliRi
rzs/jOxUtE+NDpD7e5LZC9s6YJqp3mAqX8mL3rlEsRNIIry+/jvp7W1LpJpKzvId
Y4W86sNfCNlEU8P/Y4jIZroRmzbi+XAgYLOC70aoNeKwwsAsN+FfqG2IZlNl6td6
u7TP0cbR9d/W/UCeK/f0f3XeZ+cwT0itzJhPW/YAwJ5GNTJfVrtMMuqbJW/cY5QT
uSEbmQ+my1diWh7/cDQcfEZuvvEXyxLcLrjJFZZHNrqJUG7D4aDOVj6omxfPRxma
5Q6i/P26OkRWUx3ZUjC27de4O0Jwpx4lSsfW/dIEveQFDP1BdW/sFusDk5eFhqc6
ADjYkCSRhTFhIGvV0tnYEtwEfpqb80QKzHRLS/rl82rLpo0bpH3r6lOhyq8X1Oez
3gium287sLTmMOise2L0zkm65dixaJA/dqO+MKoiu8MVUiYj0vt6cUholLbiilaZ
U8MWY2VC6cEzEOkvyW8c1EpcCMPN5+73Vff8uzWGbHnry3eQiBmBwi40kK/0UaXH
FBuc0NnIbgOztVdwTXsYDE7MucV18IsTJRiCRoJUP0sYG2MjWeGRJXMeLVeiQ8fG
TJoopSPRjDD3cpM8T0PQZEijAQ7PqvPO1fDRhkC4yKHmd5u8EHzbD6fLMCzIfeNK
m3qf16O0SbtslCVT1I6IueRt9ak7QskYH4c9TQGjXXEadZCeXT7WsnVXAQhAYOx0
sffAAUCNFkmqbfnZENGmkK3TId8WEQXeeGz4Xposu0rkfye4Zq5x7KHv1TAC2gEb
DN6rYu5N4fN17wvMXTdhdphBXygu/YtfRXIkhs6oIHywurtgqUxY/gzvtuvBKvBN
sjo8wXglAky7QnMQ7Ym/QsuPoISlmEDKWERLJdSdpxpITXoFu7dejjAEB3htS2yw
ZkXfOpxDAbtMrjJpy67jTjm3gP9aQLIhBpIk591vJYZBdLQ7LxLzdb6EKnddkG4O
Bd8j2a0LGIcXQ119Mq9QlcR+KrB6XIJ5v07T3mJgyPSVMVazHTGcEqszvWX3+en9
k1cJa/4GG5gWlErDP4r+cWDWAHG+XW/P83hcH6GYyeDv0hPxNlMJqEgG3KMvzdOj
Y1c39+eXiGixjH8PIBLlyPlys3weicBw+nRjH8UL26GUVpQbbh+jz0276UYeQ7td
I6+DRvUsOdRQ3vtEk3hP7LzpGml8bP0XeuEXoAGN5q8k9sSYViHAHNLy6UvUMv2V
5lx6tcJKYDbrND5xp5rtS5vbkZ7PzglATddSqD0nbhzFtB4f5UG3cl86vxoIYpmH
/7SP5nzHRFxzZztqbSn2m0ajTnK97JR7mUQ9DnmLk9BLAThgy1ukOSvl/iLb16hH
ogg8uvQqR7wtSPuPGh9kXiqBGeDtyAUTHVGCqO5kqKxVGqUVOSIJJLUmA74kuNlx
zw4diHIlE1j2HA93Y9msJy4JRs4rQPGSkZGid+pu9GsmEvRKK2wIT2gtTcdObrYI
i71KxVioPc6httJePZu16u9YeOzBISiLZcn+tszlyv8KME3BvbF3SB+m7n5saQjP
TmEVfbRySHR+ccz32/ge8fcmH01b5JWzAGPqpldaTNP45lh1GL9ClunDF8T0gr9z
mex6igSwafgm0SSvqghxEOV4guw/CcaIHi4KlrHuqCGZiK+5uvA9Uq7B8zUI17/p
czT2w9/wzm+MK5P0nNrmFNF5iSVwVIfPd1x8XaNcwdJ5t3/buf0HQOR7yiwecamr
aurn8CBOSBhELJ/tbXs40Ku+YOVAuuwDAbFu/Hb35qT0icbYgmaSUJMZBlyd3/hL
bHJBPB4TbDBFd/H1zcMrJY11EknhiPndjc0uzZCIlLhN+7HtYrbeQfy95fzKS2eK
jpOIFiBJiM5CNRKsgJw95FvM860xrJ730E63NBPfAqapJ7uamUcY10ctLhyOXxZo
kM90gnHO9v2ADjSI5GNJDQFvTWv1YtS1nk73sp7PmL2mfJbIdAjN1FmFhTfPsjJJ
6CqTPPdc4tQtfXA1KlewEIcKxaTxEIOTJdxARhu6ftyr8HdPUFsiK1MpxpZcOmNf
CCWHqaRyE1wcLjbYOGyACYC63Q+mV89OxKTpFU+Z/hpgH4qnlMmOd6ToKFSs/hpf
e9bEGydjD/e8ArajjS7GLixKRQ39wLKbl6nsBlfHJD9E+gcuBPONVF7Q5sZyQkZF
UoQf/Lte4ujsjumAZ8fILr0wOKwn7XX9mdsX3S7i6RODnu/PwVsL08/lZ9aODkd0
HrUp4nGyefZCWN1Z07nQOLRleww/HdDalID21BZ/V8Zt8cDUiASdIgjpQ5k+ACNW
6Ar+mNZd04WHr6vtcKM0sCq079rXVSYDu6gC4cIOaDpKo/P8K7p2+75GKhxk7Q3P
g1hKUlni/IAATz+e8yRBxFE43ZvLle3zdOGKP/94zQVkqxpCgPkDA0SEgX3ghYpD
J23bjKtXdxHBMooqDC9/5Q4T10PNAqy31pWtiZULprxdCMl+VRlUFDBeO0uGWWJ5
18E3JKiNs76O2k5RKuum+rm+GtsJfe7KNnbQUPjqeKp0l6oJ0AhnbwsS3Qg0K3GC
0ep++E1U0Jni48K9ZiCrMJ+7gAk2WrKvgq2+T9otZVjGgapNP6ugMJViOi7AKAPd
qIkgUifOMx2v1Bwjwd+6cs7CE2yPIZWTdDwBpMaPa//wbIe7x1nUL817X7AU6uIr
eZ2CI32wSPmFLIcTKx1cV2niUpi1bSALSo00xKr1G040r+ajfNE/shIZC7DQQO+6
jNM7yrS6vdhEapzASBNGXepzhoS7+YR3l6lRCrBZklGMBKInNurLMXBdDKnEtsgj
0pMxI1PSfRSklm+xfqxHNgVc8YlJw+U+1+R4wNbtwLMeaQZSJbnSjl8HCMZpSwDO
A6KWOD1ZLQv6D72a1+Qbmnz/8rFGTiUDXKhLCBOkhbHRX/mYcL3Iapoc8D/Ne8Vb
pa7PEpQx6zuiAdZdCKy9EuUaPrdbErR6k4KgJqGxQ3f22MJB1q9KB/jhCVhJZs0Z
ZFPupvyPoTUlIPiSyde3Nbwv6zql0pnn5aTLATeLMzK15Q/0zD5nAfGAMk5oKrDA
2/wMuNpZ1nMtx2m+x7EFwaih3bcLY+uSBuMccwckgBslJBpRY2Ebte0xw7PcqO0s
rmCCsZdxItDXXJEMSvYPKFTtqfkrTS2uTsr3V6HVlp+KMDmgfZRn0QkxqO70MLFi
o1gKPgFj50C8wD49b6Mp7YOkSDjZMIhLaJHVbCug+9x7Vq14kkQp1jsXVDaYG0VI
VFC5WAGHaZxcM+aB+f/zJ5QdnbTVRVyW/j2JWUYyVHs/TYQp7C2zihDN3vOk9z5E
jES3z+JL7efOxkrPAkQBUoIT0WkdyNaueuhTjzMrUTxzVPJqcOY5uAfsa/klsH4k
MhKcLz+Soek7eRterRhHa6AhOSvwtzYz6Yb+nywvzJHhSUIFICXxwGhbajSUu/rB
iEo3kdybrq9pmegCaMCYxt5sUojPx8/iG5qw/wvW6TFlddJGG2PEiX7muEzQdcQc
gcsSUzHZe7dWihW3D06UUOEA/5ThXSUDrjOrtR0/n/QxvoVP2G0VPAWzjvVUJ17c
jmB6y+R2sk3ScjVH1phPQnPsmJu1LQ2MkaB8cLfwLnLy6z7xYfS2KPO9GH32llfR
5bWtZCFqgtHnVtWAfXt++QVbEAH5W4qLPBjNBHc0c0jND6z54FKHKTd5+EeGwwLu
BrmMJU59MDKMp33mbPOyXa1mXKBNAiucT+sBu+Fimhyq9phKLmKuuP16WJp3nW2o
J5bKgXILuM3AO75Yy8wE5OIYyp8QB5IZCFFHWKrd7OWKyNU7/eniNRZoxyInoeu5
yyDkj948BRlcF3NpcK+Erwq3BRvf0ACrDPPFWKXOkh4FMnyik8g2YpSGPXOMtV6W
gm/zVfF9yuh3o5GNNGSGa6SNeWPybNAmHgY8jgV4X7ZGfKXKazPfCK/bvm3LH3Yn
4AS8ZgI+iUEWfl5+Uyo+XCut4yrh0UgoXQsNNXDzYHISV98Z5NppYJMjRwH6AFhM
ANN7j1JcwyBC0f3/LZsFl1Ltz+4rXtPJjMG6jTBnGg80C/7YFIWtPx7Xdvktap03
jpZUHstNjukFKrHByvOT4r1p8ajhjmwjaGnDeT2UL2dl9VXde2ZDxiWoU+z+5BQQ
F6Aa7ja7NvjFsWGitIbVtED1inswkBFOilBXJQNL2K/MwXfw81XNQbTAQF80NTtd
1Mnuqf+u0X/+Qk57UuvxaU/1M9rBJPLv4T3dFf1GaTI2Ae/Sl4BoCoyZzrb/25H8
p0GY9+ZwIefNGdcaF9Ii1bBfA1PsPWaZDxpimzfbB3kNYWn46Po0xJegYW16UL1Q
UV+P7vNAYLvAi5IK9Awdi94A1z0qH5FWqVEZdeyO/rvL3Kxa2KPTd/kE91rk3wcr
HiqhpAQoUbzqM4NTuwxLPTNZIGLUSfgC822pLVoHD4KDnhAIL8jwJZK1EN6ysxDw
+/YISvCUUj2FjxTE2COcV0ol5z9hFDQTkz+cDQLUIHP5ggEiHDrCLCC1kB4gJ9XG
ho+gGX4lAHvgc2lZIS4AiXywwOk57gYVwtWEJE2Sd3l0yHzMbUhs4VnapBHqvlWU
XwMSTlftndaZLS0AE31XA/NOVI/zf08odNwuWOzFQHisD2ZA1kA4RdxqjK5wJq1O
4nNzUgqBhm5eBshN6Rc6JFFquT2ilA/zoD+bNYAha7ucJmkzUaZIbJ/pMCVcMX5V
cn01NqEvhn5M7hRtZ8UxJv8JxzA48y/sAyFxslDzA+foALmADVvgoGElW2b+OdYq
MJz7HICmshOL4nWfgpYpTJ021aNWxd00peaZA00rOzBuZkK/nh99xool/0bv8BK9
Vmdh9WsM5r3cqCtHucAb6YeuCEoti8gLUpeMi2c7xnoy/mrIoUwjb7vYvqwzwAPT
AzeIK6q/MlRVwLOA9Xc6fRIDElXJv1gddczot0uE8qsxeRuxqZTSVNB9iM8pjzDC
AYKIsiRenk0vcBqD9yN6pAnRIlSkFDvf/GY+F7YQVUpNIhbgHl5XrIAYFmyRqm+O
l34yaFZD0gts6TYmLEkACQAf0bcBuGyblgEuYNB572nF6LEd69z3WTBiXtVA9fj7
sPQdiQClhRLEQgC5lQEKCLu779jeFw2QjipN2LkahUwiU0+VHS9PDxkRjaLHQVNP
l+yKZBFUNIeWAPScnHg5O6m/J4BX5i+GNE7muIAo4ETxzpq5738gq4vpPclMcQe1
tUZJlxdO8sDF9J6117XmG7XDWjRk2aivWtZVKA+aN/4eD/q3T1x5n0a5yZE8DPa5
KATkHbLRlMswlAP5x8ai9Moo8exAew9dzD07tiJVtN2oNXKZlzpkkiWurP/dzLa5
BB3cZIosyWLHmhJeva8Mfwbra/R36rMa7yqstE8TZ39y4CTQl7US92DtnJr/lURV
7uRSB1RsA08xQjCbjwca9ZpMw9Is6W+Lk47LWF4JT01qDwhRqdVYnQuxp8kOm/Fj
KNb7hkD+VDch9BX4JlMxDMBDrwqmNEspV7kd4U/3TYjl+Bq1XJlEG/9xf0iRxhZa
MmG1i8WOGUs35AzlNN+4eppxl72a9FyJI451FfPnKkYvqMWCE8ndRVUG7QtuyiCI
2RpQxokp4thr1S8gtTpzaOyK3aTzjyYyJNPfGlsvkkL+v0foVYth+betqnjKpvqs
jRyeu0UsJPLtD3RoPrxEEx/463A7WIc0QwQ8QBFYPjxjecefz7uaCKLDTSuUahNx
2mwn3VWqx2trQG7xIXtMqLNiH508ByHvJG/ZzNLvovh8mgjOWM3fUqlUg8ZGvRLK
2mhTcincEwL0LQgT7U8zgAp8rNOI3Bjk4ORLLv8F0qQpm+7C/tF2MyEWTAM30RmA
7WgIOIiWUS5yTPRFZWjzIzspW2nqnbyeZ59q7F2Xzz+Y3b/I90Ax03rkhRzZipIm
vlL5X8+Pf2RBA8G2Qp/e7VfNr7+jOK954guCWQRbQpyRyIYqduXpbckQjXW62RVD
ZA0Yk5XA62kv0wlPg6+RU8+iaEme4OpVJ1zRpgxUXYau8szDNI4vH8ZSBlhnK2Nk
YchtHxu7QFJIRqoMMMINVXidw+1Caw8J9IUh+d0si5h4tLVRrB4vMKp5w5CBoFPX
tWJeCo6hQ82rFIfZj9PFF8PvVsZJdtHlSBYeH623m/d9raoWqQu3+t3S4huxwHEw
OEduKUGkJ/oWIKG1gfc5n15aqjIoRkBNot4oneN2uv7hSENQ9cJ3IshKM8dEr9/D
bTDYwh6qP2M5kqU6QWdmvKmoLuRauq0fXT9ddVobH/hBQgdZE7hMXZZXZDMGLj7y
ACwGxcBKCzsXMoc/MuifrWPrwb6cX3qf9UN75Bh6alG3cVn8bQR2j2fZFG9uxQ2K
Qk6E6FxLxUPT/xJe1DMpWJOiZ6nvwE3uD6NVYdqpPaeNH21VZKG4YxfUaz2dJaBj
IHK/UU0QEC6JWw55taXULj44Tqj3lvQdR4T7YV1sy3jeOgYRSqq19xu8nUpgsD26
gAN06WspCYiNOvySS0LMT5YRQD+gPGKomXLyCFBm6zuClG3nY2sUKkbMdO5YDnMj
8pGhoq7SbRRoo7mBE4TqG1NmOgPJP6UXxuME399PnPveGBUlU6W8/DBTpqb5JF30
9C7/SpuD2To+OqDcY6um8kkrU3eiPzmsRHEsklSlWyab2Bxz1AzQJEiWO98Nw399
0xiNt55qI2MZWXMc7nvPYpwLu3/EmtHXTgrue16eE9y9lYSa+Gpi6WJwTrh6sL4n
TiRgspMoXRMEJin4UHwBoAuf4YzyrFjfYZ+a/868NPuuutcGdqIcRfpIeznNZtMo
3bgitPmzhjrnh6uWXttPPJkBqoi4ckHxrdnkxV8ijIG8STl2ygwSLUbWGZX7ptYo
/+N9VO5Te/A5sdPKZLezLepXpte3LgqMNYeMnR3nqTNMsqCEvg7p7tMaRXWRLKak
lD+x3eVw4u6VGhp7PFk0q8NjSxf4acWf2spnP6PMb83v29x8HKuKLxwr+7iWAgGJ
BF2MEeKYp2ihIDKpX06Fc64xETizSMHvgNy15kK4actNU5NGbEgGUE/fbhjq8jik
vFTRT5P4MZ633A/4EN/9thWX2l+xgvjc6Aam2tU+ovP4+ua+aCwr6mcphqn7M+RJ
z6kR5a0L9/qrt1L9w8ApqSCvDWwwLBDIfnjPpt36tZD0h4BQebIz1tO1r9wGjtKQ
a6bi96peoQkxKwGfaLmIjcqKwiR9AmVPk206/vJGh3JA3u677YUqKQv7oviol5nJ
ywRNPLxJBpXTgz6FaSy0zrK6b+pOLvV5NE+k6bGiGZHqxqmfy6421sJgbGhvRAQj
YleuFr44lhUYdbqDRYE+WrUmuNMbcRv+Aif1+y0SQBKLu+nC9T58jG6iDvEJklBb
ilb/i6aYnnF7fB2H91u7ZJht19RHF1c7sw8Sw3e+CpCruCBYVnvMqx5K4flKAgL4
zG2JR0cafQC3IwtVZxWQOURsyMtZyzNsptgeUGmCizc7h+RezN1Yh41f3idf1C7X
9P8hpJ0O9JdnBAqUcjrENlXPT0wxry51ne9YrlD7JxVEkTk0b2XovtaVJncixvQZ
ZEGKR+pISZdBs0cmFCMMPVeGkid5ycILSSnJWTT1ZaWZzkrDwITh1B4ZzBvioJPc
++tpoegHAErsOF3lxeEragHvBuKfoY82Eq2BYQNup3gT1Tkw/cPoxx1dTfO7DlQ7
/jwyKBbv3kFfpk5Za8ZRNSMSPyakgYScYhZPMkcjv61ETmudWFUaHaRimbVmLn6J
Uczva5BP+xYGsHoLI7i31ROXqFNofxJKHGcKkPCcQfQBElpZ+UhaNLe12jt598Nk
7yKl13PIjdam4ANeVWoA5A8Rxgus5MSTp4/c94/ZV37iiZoglu+Saj1Y5CCkDAF3
UWgrDvWM2hNSmNtJSRWGelAfhsD2yIlaXKt6RNYu0jSnETJH8RfUlW9/AVEfFr5c
Qxbq3nPnCwp9O4RH5+WG4wY7yOviYpRvMichy1zoTSX43vfIbwgvFo6LVNmVZaNY
YCyE5GDAzplJOj7Az//vYuYMvRdYO8GEAvB/k5OHXF6pf5rTs72Qq10tqz1pPLQo
5rRTUrba+RsPLpw6uit2yASFeYYj5AR5S4+FR8Rb3qBkuAKaZET0NgZFJpW9UGsv
LeY3KgYCw8oXMB/kUEkC7aEncgCYC7Da/XQpkjWzXNCdJfTlbOF6wIUOJVKQl4Uz
2NDkWqLErfsY5fKsaIXaWxRFzs1UzwRwPcexdiAhFwzRNFiv7UuKpGsD29qZ8bIQ
2NGdWeikwMc1wU0yOYTLYO1r5Fsx0X0c8kDZUi0MLLeETkbxf1knYkxkEeYDo8hV
0lrW9KfDn6qJiph+dbGwsBbJE9PQF1zCdgGAY2kiaLLYx0r0z/Jrby0LX6CCKTWx
BUWXSLm/PKht8dDmsX75MAHNZsEL9J1qsWQwy9xbUXz9rS+OMVgK2PbbSJOs8k65
tUmoUxu8KS5IfCQzlB4LQFWW1cooxTWUgGI2AszelNagRzBDKZ08maYmrXAAC7hr
PQbpN4kgSURkc7nw/Aw4a8Y9LmS5E4xc+PiwurXo20vel1cUzImYO1iirsfKvBFr
nr92G4n5+cAnLw4wGvbiqizyrM3h5/leV5kYNM9nwSXzGBURwzYGmOkEiQt6bnm1
F9n6X0+p8fL1XTO9g95i0ZDVVpsTkyE2OwCniw+BSpLvmQm79jJBcwxyHe+ZTFuN
tnWVB/QGn+XUGu0dUvanRgCohuuHLNKS8GHa7J+ULHLSW2T1Y9AXd8YY/6pjWKpp
8AIkPQlDbR65dfNWs85vBTWeCZF7RBY+5yAWkNOD8OOeqGu5n5gXDpL56qYumvi2
QQty8zoibP1Og0MjPugoX+Vw5FeceuMHEjyvcbhev3G2YrMXwQXZtBB1N4Zvoy2i
PF8+tw6ZmODpH+Ez2ltiUziyimgdR92rn8M57R3tD7qp/JEh+oTWCpkBo/DjRM6x
mx5vm80AjBU1ymSp4ytxSMK9fT+5AjIdMHpmB3dprkK9pVYDjuKCEEwjSeFgZ7EK
7PiDT+kHcXI+AHPW0dSl7Srn3tqSVOQXhNC27nq6YEEE0hzNgqFfwU5ishWsfgyQ
YyufYPTMv1/SaM7wyzVpvez79RCVspdCd8zVlTFNDZVlNEvbCzIKXISNrVnONLms
Yud9rlOu6+kyiHgs4d56mXS3fWWuiru9y4Qbmo91C3e54Jpu987KtUQxeYLDD8Cl
0V6bF1xsGBGl39b3oFqKA/x0uFcv3h6Ap9Yf8L9aKQxAit9q3Khx4vOMjXQT89Ug
1AgT086Ev5nsM8pl2Gz169aUUba9OHsKl0lUhhSe4dpGi2v/F978auHn6c+M3ghA
BrmZycxH3/xNMqJLCjRhTMkIjOmYmfS/vJR92l2XUwxJedSI0pyBycvTgPx5dza5
XUBmfNg1JHeUol7I1s1bhTjjjzFyIK6YTylpiKosS3j3DXp41qeUgwx/U8YPj9t9
ao7NzeXHzLyoW9hBnlsBM3EAwAYc3dyEaZyO4+10hexzWlZcTWLX07kq65ZGQWmv
Umwm3C/+DLluKuzmZdovLrdgS2S8yc9lw2m5rkITFcMMtuwcF1sicDWzRyJeRXQe
rGZ1CTcGHmWRe+kv76pIy5r5lGaEl57vSUFpOkf3bhjBPd94IYJGVTJZ21Cp42f6
NP4DzwA/Lb2b1lBJS6/lUPKS3C90VIXwxsncWxCnf8VLiWBQiMgTHwQ9CzVNqYR0
T45FLNCRI75dZm4uwkR7SHDqfHYwhiD3JLeQWJB/bvcfze8oiZzTXspjQweay36W
7VQuvGiEZoinJCkmZ3o8bnlqyG9xn+x30AmPL/sXauA6T6VFbcxZ5YG1HDaQLCEq
cOwRxaHrxD4jsEqsss0CCDt0l9up9a3XKH0O8gwYdzV9ErlEg6Z513wE21NXJVHn
ARjAq0yx12awvTrEcLJGnXWqFL71pAIm1LJfMvT/Y+DwKJ/il0LVZKCdc8BUHfRq
vR7QxToiAG1H359srCqskms3BXksp5mR3ozCZDzVmHDDWa7uAkNfXVSBTrSiGYFA
QqV7vfYBSkwJjtmb9enIfgZSAAy/wLpOB6cx5VZVeghDbV8oOF1Fh9U4jdPoYYqs
nSDOQkzs5L8+4L1pZR5JPE3QELOljvvuC3EWl9oqxcecNQciL59x13lZ+tDhDFfH
JI8MpEQGvBzTCofqqauSbLdCBdtQfRktMzkGY02wk0yHFX8eVMJWsiIn55fNxQN0
pIB226nJBhMO+mmduPqaIauMvUzuYqcBDtuqSHvL1qtnqDiHAuljCoh0n7foVDHK
vyOjl+5ZBba5h1AdLPUeoaGTonXOzHQeUjaG8ykQacL0q2KmqYn/T0Tsewa6Lb33
0EDdj9wY1SXOhykvbb0RGMZwRR2Gty5ru9QOFvQLK85KyJeu8o0VosOiQZ1JlF7i
OWsduNlsILIIkU/mSSbpWE5dJbRtvhmVuhhhEH8IMp6kCuwRAUHNVjtarSu9oUpI
/vLrctjy3OmXP5bjfZWqCRUEtvhRzpp35MWSFKkGufSYA6A96bUlKxXRmf0SbG6q
dGp6lT7K2l5MwKSlCqTPc+J+aX4mu0ucs7ShpTFvtJNqBeJRhGEmQN2RhLOASEkk
R01Ivfq59DIhAl1x+vv7Evd0+8qFKaYmO9P1wSV0IfO/SRnczIjlf0qlTjXvCJyA
jBIpyCjYseFRPwPZynvZ1vOGQFo2xMq9XrrVz4DU9mCvjJVmOEnX8IWnbP8mcEXJ
MLJuuUtCPW7zkoucUofH2VES1MY1bt7E8wHZwCb6kJ7XjY9rawWi+h22LkvEqNwL
eqBNUto7vI2HPQICRzbb00v9G8rTepgyOOOyTCthTX47guzGwrkTTrZB6APoDa1d
FUFY7YfuXRYOGxM35XUs+Hk4ULNEbFlEVZT8JwEcthm5r66wm08QmtNci9FaHUja
r9NQPCeyHGSNIWSv4nyp5K6fAKy3lTTUO2lp2khC60Ud3ec6I/Vgo75AxwCzF35G
Csk6uw5A7VJzlVZ9ri6lwFWzCupYsqll1iRPJSXFIHyLn++yHButpqoopsWYl2aW
fkmWXKZ13FVVrPvQ99mxCmIl7klOQtCcoR+rpjjo67kuwsGKG2BROpK7Eopf9R4X
SrvFPrEj7HbC5in+LbU9wWxPoYG8ImXMnHepuI90jXduyirs4fatLYoUQIPIxqCo
OkNcP4tQ36jGSOa+JRAh9qtXDVsgyP+umc+tM8KJQa7dt5sCYHdhRDAQETn5Xrgc
q9mSGKpsPP+m/NS/AE+BYRPM/1GInSDNHgZYkrFSp9/LQq+6EP09u/B4AGCPvFoz
VLOTQzIqLWy6u1rus8990Umkigp7BDn0mrOHfVaANLG75nI15Wr0NZKbGopmMO90
R3KPVs3ScUfmdRaYXUaQJ2IF8pc7KrHYNgWiV8rXJwnc+fW8xXE2J1LGk9DiZ4Bx
4VLoJ9lSG3Y82WYN4cSH7tWBsyu1J1bQx0Ol8I30nGdsnQnAER7T+pVPQZ6uXUdx
9lPBZ2gE3m4jT43EXzKTvYvixQ3MYF1EPKTpa24zVcsi4ooHuCuSAvmLlAnAvEVv
PTE0tlCpch70isU+XY1rMh85XY/PZlQcD7PwC9f0mEWMiOE7hUVF/fCHXtdTKbz3
oWBZmuqIWAnhUFApn5Y1yogIxvJcfD0kbwtknEEA97TAeYsTq2oPwuR1Hl+6j8+C
0BP8bS+XgAtWdTmeNKSxoeUTT5MZ7J/AYcc572biH/UEQ8YC0yWlatO6VgXP/Oq5
rt4dnoJI910H+BpByzs6SmqWfffxcGlq9RKX5I9MwR2OLAY3v3obW7hPSfrr0HZw
rBm9h92DV93uy6JXlQXuchPC6I+d63/n8RKOZPi3aTmOFkKMPhg7NAV4hmdKJ4vi
BiLGS0gfxkUUCgsHLhLVDDiZ6FedNbJGfsIJzI6LXvp2T8y+G4YC2IvvA8zJUzpn
2hdTNHfEbkyTu7+peWZkOxlcxoZzMgaRg+/+B39IR+BItk1qCpHuxgevXlx1TIlJ
EOfbBQZCM3evoNWahnf0iu54OGbEX2qqpO40v1oUPSurX4AukdxV684hqxa4cGCi
YnpaV7j2Eo08E80WwrzonrDuOVFgYFUHRYMVnVLyN66K8pMBMAb/h2R5HFqOuHuf
HAvXHYw0/qLQVWiNph0ejCwK1tYvvn5BkckCCqf47qVgzH8f8t6S+7OJsRT6gs33
e+9eF0a0wg9WDlsRIW1wM6jXVFHUyS+Px/8G7gOOyyArgXzoQAcP7pkt615L5IYA
QS3GNR9Ol5MDPdm3mvrCQu8fTnOHbNtJRhRYlPplI1JQLQ+E9gK0jGtKN3iCh3LD
GaRKgweT8ZejRdorEloGDyizDRRn22a/B0w3s84oVwNFk9IMAV4YyiejcDUmWJ4Y
3gj4E2xycxW7usUeCKWKCZAbKJwVZcXfdCneVMQn2hVItOWThXNpwYbfI7xCwLQJ
O0eMiG42KGV7mVvNMx/V1M3eAInXokdEhDtz8lnD0GucN/qGyH1wy8cFKnbQvXcd
YKY00FKFTtDAWA4a+jJFHfIPsYwjNppizgYV3wATQ05GZuDYk+9jlpLssIYHX/xs
prOBIXGDXQ+CXHO+MwiiLwqLF5EVK4fum4B+EdwRU16fAQxkZuX4gRn5Mz4Fqz4z
7kM1J6MrWrcwJivdwYUlqdFud9A7sn2IHyIcwtK3uLE9z9+VCIw6LxFspsIevzLu
jxHmqqm6HBC5qCEbJfQX1IPpbShgtfVID/05p+MMeEM5g8pg1k1ZK53Ad+QZ7IDg
z2JO1IFcjIzJhxu8mVX75dcVpbK8hePLe+/U8Tj4spWHvYKn3PzPNOnhKuesB/sv
jX4S6JML30MuC4NN3Nf3gp67oYasIRLe/FtJna1PgH2mV1sVB7hXIZX+ntUpPSKM
74mGh8d39S3xqRzuIf7fqsMfJ3DOwEwi+HLhQQw+9xiVOE8Ca/UDWgoLPPSwBQKe
UVkkjwXaAA9HEhwvOMOKpHvnKl+sAJ47LckntmqlXhSgN2M6V8FrvrhoMzsfhynk
7vChSEKRN7PZE5aO9aJez3eAIvDwmD9VymzHKQTZHAjPflKdDxMbvnGt5hwwIlpw
3Zs7w+PON8jZAE9ASDTnbISvlxRcNIEoeytNo188qATItX5NSpQtepibrColK0aK
t32DPPf+IWY6iomC2Gi2ztyz6zbqnZbhPUT1NnHBwRZkKxzJ2rqj1NTfXVt9tKNM
9eCNn+SfVEMVkvK0DjUL7w5ZTLX4U1vjzOx5p7cY3cUC4KQs32/L5YkGVyEwwd+R
QHGuYEefDfpI4xUpyXm/hFBexdlPOE9wxCftijzbR6MPczu2q4OH+pRVaHUmBimo
hzvg4mLaBFgtF7TnTGdRHPfsTQBo9YFyNYsgTsjjW9SGmiTktjlqQXse7L5Fw1bh
kD/4TbJa3PV/KhYJgGJpNwy5D1kfaR6szFLqX9I/EbXvd1GexwFkEaeYifdubE4H
ipRaXnfQYxZZ7chISClHnYuK27Jco0is32WQrsDYTSLAtOU6gJ3NM+/l6zLEl786
rPfSHQn0zSplAMDOtzBw5R6jQnvd8bXLPu69nCt+PDX+Uuj8OJb/QoW6LovicA0U
OtokcpP/NTAZN0oa1kupfMsF2kdXW0y2ccqaaonUSLDBK/6UrOVoWRJsygrYpeeb
tzmy+5+Q1U+1FMuGllxWdRt77pc3y7oTCTdww648osCwHohRzZpruCQtWXtUCSO+
K+FBuBrUJSLXHzQIipc+BaHgzyuHdgD+dkQwA9M9+fnXPi5yz+NfOP6arfPxtWCf
q3XmTQXtFFNR9+mQphaZamR3AAodrXdOc1Md4PrLu+7VJhzE9E1+yN6qneXrL5Iq
/mdkb13FGOhEgZ5T4ct43in5S+5fmyvxdackXABwMPaO+zd+391d9wArhe8KYDHd
8YW1wHLdVoDABqluY80GTxQlFZ3h33M3LsExI/4rPurst1hubr7YXWQw8S64kbDM
vRsOEs5bGecAK5FXZpWwVB+qEMbGrcY+MlmBGTDdpt79rP4X1YH33gq97h8dMJpl
sOqZCtFeAG1TajTyT4gWJL8V3Wsk+IfT2rtCLKefkJjrtzSAgAmMM9D8nCwLv0qN
xyZnluiCVUGnnJZYsfIMIcF6xLnKwZi1a3IXJ/uGOs7r4/7JuNPhgcrzmxL+hCBO
FV52pNjaIUdPXwYh1oUiXk402Q58euJ2GoZbBfjMF5Kro1GyRBVcFmt6n6o19HVl
CyoajZjQj1Zi6FqfqxYAuQKnp/9m3gMT0nNNkxIZ14g5b4FlpB3BDamv4O7P8fVo
O5xeY88MstlYPuMzh8tai+aqv/h0ZhySXieOJJLjnGMnZ/Fy6FDfaM69usyqKSoA
b1HGpqAgmNTO865LFrvI8HjUJQOsPCS283bq0uvAF7uhBlWfwDQD/ZDF4ACQ/Cme
LShwvF00NGCCeVgy193Ea16tolQYaJAs/d/b3YXbAxhfgGP48bsgdNV7jRTm/Zlj
xUWASDQqb1C31sM5ZnzlMQBdaVesGgHZvC7E84BQuMZ0uWKLpaFv8e79/JZ8cfP/
KtbL6JPK+kqCp6ZHTMYspgVZAkg6FtqDuVr6FRUrlCw9QD7kWZQANxvtaPP/DE2s
RfYhnXzHX4P+2O5BNXQtgPwxPApbRbfzhgpciU+TonJZoTHt2bpNLWnKi6P4v1nY
cDq7k7AHjhW7+uNdPhC6kX7hrVtZgZacLLOF/ACpa+Z3646VsVcK0MkBirOg/m3s
hG7A2x5dGCbvBnaXuA5k8TF87QvBKDVlOZ4jssSBk4qNI9KYkUvV3N27fHmlj6PL
ZhPAva6+kvevXDbRtBYyILaBKf7CQ1pl9wAYbORcO8/pj7ev0zo82+XMKMnW6prl
P+z65wmSAGEf9jKEcHC4Fl/bgmqMYUvwAuYkejwOkfcKqN8N4I+1AfCI1hCxPmKj
kkPjXr6vfxt6gH9J7C7fAMZynABkM9m2KB27+2QFoKrxowTQM37JSJ9LNzB0Ntbl
fhbSiN/bkV7jRyB4Eost4JbXIg3NEyCqHocW4FRUTG2MO8JHC5OyR+n0iXSBuAyE
X+B2fx4V7/QtfnLAsBchkFX0eOABKnKjiGn17vXKUEiUPvQvZXF5ecSptdztRAY5
mxrkpEkff10e7iTPBhcwCyWB1KrsNBcUIutjXPjlKZ4azcvW8AgZw4wrspDI/KVF
NL3UyGtXmggarEiWc/nS41RvRNUiWxx8NHlzQypioC6FgXNs/ottqqje4AQEvb2m
8UAee1TKNpXO5DhWui5nH3Rd6UHSuINOdNog9RabaZ+yQXLHPpHoCQA8o4Tq6LSb
yArFuVZz+1lJk5iEqYSaCxO4jaD5Do5KCgaNPKq47VUqjERMu4dFWdmQTZtWUoe7
1KuSFOP4dOZCx7wIlte0MSdv6MMioRZOxkhWghFKzVq6UwPnEN77UQHKaQdIE3A0
acStKI6Bkro8JVk9XQCNRy2WKrOuBI+cd8G9chmfffesKLg1OloonuAp3cQMRYqy
68E4yzMmf9UbjhGj9KUroUPftsbq7NcfRc3J+o8FzlU+nZACo5Ten6NJyJVsNycJ
rpyywK2mmNiMpT54eJ4nTT3FTZHrJrPPwvC/+NZmFvgskmrULJJZ5k/Q4UAu5u8L
sYVug0s5ywspUQbu0iKp4Fl3RX6/Q21RVAk/u760SZElbuo/QbHHFHHD/wdlN/7P
9JT8etl2H5BuUhYLS0nOorYhb90C3QDFqmClnNYchkot1OvuCitaQ9TiLxf6i23B
iwlo7v9Xu/kakZczFCdsT9X5eC72AQziMjK6LFDf7U+nA+5uwLHoTfFa8jtZt4gK
3cxQ/4KjqsCOMugRY3mnrVLM2w3/RugKRA8ghwFWZYJVqlOWbq3m1lkehXG5YwuP
WALwpRy+wJVW5ISJPnNLR/4rQmilfLgnxdaGIOdjjs0R6YYvahLoTHWhOpu06i+G
6p/522jYUF75+vC7uF1nkFDImvTjYJa2T81DdToE+dOQKWQSMeF9MdZ7QuL8WCd0
8cfJ/LftLoNirPjG0RdfdD3Jyr7b4FKG+MLWwG2VGisTus61VbSAY/7vjo/168aP
It1pgYMJYqgFuQYBDE4X2ARsbULBQBUV/HI5Sr1maYczZRn+Aqny+b9o11N7KZQL
9hfMQ0x8ysI6ZaNAfOilkPViLFqWpELOK1tPu+25Vkf6yrDA7t+0mr6ObXtxmxkh
HjVU6Nd/widHRBiVmKahPW3lxSiNu8gu4TIeZxOBOaaDixtkFuMgtQJz4IZEissc
Y6Yi6662hOdVTBNnRyx9YGuT9MEBlISbxT+fcVxk2kqQZbUEt14OPZ6OFbODsoqo
yAKOv7PFgduCyrcj9Ij5y+qKTHsH6fMv1Nk1OlZjvkFxGxnPIIIYdsALm9+jb4w9
BOtYxfco28YQCLOY9RIvBc9uMJMNWr/m8czQlFFmjDwsorOGfoQao9W0LMIFy94o
8gDHohDxy5vzqYWiTBXOHixIQlakFElrXT+iEP/Sz8fT57E3nJWQAig8zXhQHMhJ
+dfN/7bAyMCcRw6wMsR40bsJ/PiFfoVOSQJ4ELt8cxdFiAzOYPviDUlnxV0bDgT9
FTN/T3qR3Oz9oYHyS4w7MEglDu2snPcpxyTFlu7zyVSRYJZBTUWtfkC9BQSmTQzx
HL8Lyl6mzdpMtS/Bkv5Zfgr06zGZW2trGigx97aYV+YcrE8SUgLk0V4/Tig9E7ms
gOjy3AQK96EHKVn8WUdLd4u7Z/r0Ph6G9w3kzSkFTphm6ZpT0UPZPzwYhN/8+bMV
2NCv8vsZU7coBK41tuHnJzClC5f44FZJAQmaxOHnicQIKTr6AuFtL9qnQ41Wne4o
4tiOIFD65WDy9A2I1/unYaXdZy0q0bXej2I92F0Ro9rUJD6EIryIFzAOXXQs4pN/
qo01nFf1SQgaElF+zBut+6GikuVtXBjkt8aRJDv7fa6pV6ZcULBktvBIDVBet4H9
SoN3SMXoSBPm9M3OH5g18f0z++J5VZYcMKeIqAJn2gKj9J6RjrnZB0OWHbWsqp/O
US9FuVSqeqwqx4ljloqm97qWqdX8yxl0wHyY4bnuy9LGHLmGVQdfH67cMbO+OyMW
Y3c/huP0ioG6JfXf1T9W2ZpUlMteDjRsX0VqjexsaRSc9V7Ak+AeCcF0w1/zZ5yb
lVe6OKxTVpe+EVBjdijdVVybHI9IADb7vnK4hDO8O7mIrsr43NcIk8boflTGDyCz
I1svosZ6fQ0feaGz01tODEueoqsyU5A8/yD7C7AMkxVnE1vWjMXZ0nuhzARHmbjT
Cj7ezQ9v5j5VuNMLniwCqKOh6ug2XhtDshajpElCz0qMGt4iTPhCj4ZRcmjOQl9f
klOzA+Ysaelf4vxTaBIOxYgSeR10HCkdLliLvch1iEL/Koa7ULQJkPSJqSvDHhoZ
tRO/4n99af4M/bRURT22nGHRNeY3w5y3vu1QccIZi++vyVYNP36ECHeiNChTkZzX
Yv/WDn/rjfvguH2lWsXwFt9Rdw2STRurhuBop7WweDFTwSM/GQB/Ibzp6W8RozmB
qdRmZgSxArGEOv+KsKt0a3MN+rczh6ojyHfy//b9KyvsTVsi5be4ytM298TJuZ/B
bLpHPv5ieirFeHq3bNaOIOTeufYAyLEFt0Wx1Wmtov8Wss9Hw0CYjwPtFt++8sd5
/gyCoTdMmrIzjZv/iFS1IHWwg5JL1b6ozg8O51JXWl3xpqX87sA8PV5sKAQzVhtA
475kZTgEF9BcC2T+eMeMLkv0aks1D8ZJxSipjwXzWJFpyd7lVY5l5hB6lwRcG2eB
moh4CIEmSC5N0oGdq8ou+ak3z7oLeIxSgl0tkiAqAW40oGi5/Q5CLZ3o/ZQe8UwE
DkRBUJ4floD9j2ygYH0JUv+JXORzkIBlShmrRgo390vMYhRtL3b04Ci+/95Soq2I
go+1aRXrAovGQtLK8RFJC9itcrvdUpxFAyvOsVscBzYNmvE3jofZIIsi1qk+DR+H
yK4wNasjI6h1BOgtRVrtEV4gXqENK8a3M7UHxIMpsPbUoxnR9X+Qv6GlxasOkw9T
mFCq97SwfmkLaWcZcmSXJUk12ZWvkKuhpmFrANSEHktx/FHnrjr0oGbaD7rramgV
tnsGXH+zX2zW/Wzsju2xuxOhVaAIaflOox8y+nRrZ1o6ZsZsavnlrmPfVlTbUAYG
VfScqT2pb2OmM8PPBQ63m4UTP6BJy6QjRmtNDAML7W0bmRyYW0lUuSdB0D/w2ucs
JZisRIRVMAFNeA7KfUPcKDbGSqJKReOkKkDrqFszXlyXKbXnF7ZEBCNNA3Odh+5U
w2KK5qxzzK8yehUaz2JMMU1+ZwfXRvFv34LpVirMncMkuaI8s0AnBe0nadEPc0vD
3vUokAA/6DF3G2NOMMtYoVqklXjJ44cfoHEuLt7CcchdJysaCq8eeHqWeRx47LK+
Hd9MS0BvKcD9q+lv9sYNrQMEgQ1bmfN5VhdA3+NK4mgoXyIW9YSgJyxwRqc6O4vY
0cmDSe128KcwNrxqQuclNqLCkLHYcM8mcarhsYBGw0lMbMUHanclhgyhiEl9N1ZF
IIZlJIW4DQfISBYerIxeFgkVkOpzOE/1FTNXO80vsFj2ecHjlQXyqr4zhC1Rw0/b
YGvQ7HqCbl3g8jaYiI3DLczf8p9WTqtitfHhMYXSsxrVBwdbXEyd1Wh9+BML/OHp
7am7vuWrxAHBUNPInn4qNab7pwG/+1JHy+henMe0D7uPwUizs7t0W0EVkxcVELIN
bqJDVxeZZ1RxYyzrKkEDwxbAl9Ls6qVyjdy7OML2zTBSUM7t8ECdCcag7rCkJOCN
3wY2U4JzzY+mkIk6vh9N1ZHus5Z8u6DCwqFssvoLe6iMMdGXLF/aSI/B2mNSjBHO
bWhV3q5A2TaJRyFKu3Df48Z4QM0MpcEarV2/fJGB8be0r+votIxgPrMu5YIJsAS6
Z/y1u+Djn5kcwa1YwBKsFlLM/J3fz/+HLQqB1txeN8yAfhlaQd6afACEYALvTjeN
1A+ffw9I+4GhVIG47vZlkGnusLH57PWo1G1MRDjdVIwVew0wu7fZPx0eIs29wWcK
K7wddzk4YwsL1u3fztzAbtHdsSJ49yF9jdxXHiGkGr7utQkL6Gmm9UgrWCrL96Tg
9wuV+NUKqD0L+YyvoBxqpl0wAbQjgz2vtcTk1w3AlLRRQlppFYdMW14iUVwSdQkH
Oxy+J+mAaWqYLWTzMO/rswkJtI92n5ai1OPDxOHv+qzRfrCvxd6AlrTaQDI7nNHx
0TJTXnOop4qoMbGH75/aeaYZzEkHH1if04LYlRcCzuDWNbTTKVBh9fZCmH1x7ZR6
uzkgdj4GSbY/U6jEBPL38G3QhzurCE82jZ7X2IKmwq9lv1f4yP2XE8PuSR8bMPlR
OvzbInPf4zGQ773mNi3aclmDdU19Pj5D7JzfpmLay9bOKvEztkSs2qqzmI1NGWG+
EgHvx+TPQCFAylvFRGgKLqZ0x/K8Te2176C+iPgcpBR0YJPfzlIdc674h21dJ6s9
QzAzZLIVepRJwfPCMUxyGQ5Epvxp0f1spSGB/POMuoTvX94H5XI88Dc16a9+yKEz
xEkJskAQAn1/VVExacxmWS0uacIsZClv6guFvYvqq7AR2HTINppftX1lH6BkwMKi
/25/PpT0h9F+C9u3jaAXpQLqkE8vSy7QZIc67chZz8EW6due8IVs8focFKvgbwsJ
SobiyzzBtpzwhNPnonNwNx73UX/+YyNUMBRUGciyUtKrsXIdn69Zqj/w67tYwDK2
xkXprrg5GOk4y9oyY2dWzotqoPDzgU07sAPVtPi4/nW6jp8cU6fnMufLv1h6ITKK
lNRLScCE0ChTxKjGtRWdYAEcOet8bZKLPeMFdWL663qtIAnn9qRu7j41/ss7xFIl
/SNSyKFOZm4hi4pmJEQO9SZSgeXJXW15mDp65AdrfpmI6+IPUtsOxsKjGe5IS3Kx
xp2Hks6qWtS4Fj5ob7C07i4pWhD9a7p/xWPh7UGIpEIObsdRsBAiW8JS9C9oM41C
2ku1/gE98uh1HcRJtogKSlXcV0nrx0EXNcW4nZsHej1SsjXHqAN1b98VGRcQZhrY
Qe+mPLt9XxDKSzSBDdaUqPqMhOCJ7RI52QKC3WxeWCoRXbrnXFpr9GVgwXQIGh1H
48PqXkDF8+4mbdR8plJiMryEltp5Dv5h6KtsHiRxJtk5P12dUbs1UnWj+RyQXzff
5YrK+/mMkM8f3R8tTAvOvqVPi/jDw2rcHGI8bRDi/7gbQL5rJf7xeuAjy443Zyr3
d4rU61PBRYIzm3CgOnGFsWxW5Ocyu0pNRapU7WTxRFrxlpLDgjIQz3UdN1nMibKj
N7QziHMnbL6a+REWBgQ9xkILaZkYGiWWiZxuw+Hqi/8SCoH6o2wIrfr3goC84LEh
7wl9/J3aY2qz8s8lhSL8etanLO4Z9gAKiX+wUO2vOW4utZeT5u7FC94NIDoOpG8J
2HkmUApLc1TzYWqkXH3I3vRDiqK2lhXBWJDrV9ptFTHdb1PFhxknRCaMhPsLGFSD
IRwhY2TQy5sTMwpH69oodwgJsYIFbwowtJbf/A7Mq1JTtIzmg9fty+WGIUoobUV4
udGK7IfyuQdFanpPEmHYmS0QPhuzeYdwf7tSc1r593Qt/jgkf2C3sh6nNqJWZq6I
ZLSlQSnqZFDdkOKer0VdDIVHXd77iE+cWI4R39QptbfWpGPz2owE6rr0IQ/+RVUh
PBuPFDQNfypxLvkxlXaKO7vaL2Rtfg1Bpoc0Gsr4ueqq8f6T6eBTq07KpXu9lQ9V
dhE2Mo0aja5gzpCiMQ0ykILD5hYcoeNI/ZqD8gN3ImkwahKxmfjUH6Pk07SRKAKb
FpuCVvc5etxTUo3fZpFAJUTW4wmnjX9TDgrWjksGAYwVQ4sS8oHbSsqXf+TW5yXk
oQqG3+Re+WkoIVD7dDnL/37BNpW71RCJi1SNi6u+sJxgCSFgFYTHmEF2l+OByRxi
aukVu33lcRxcqm/Mr51o0Xnpl+wLLy3qQS6TgJuyLl21nxCxRh4Agkt+GgEOwDm6
xKhEroIaAPTQeaH84FAYjIwx8E9td3LrXcLGLPOwDRkNZpUCh8QtktF+Q6pFrWbs
k2CEVrmFgZQl3bXxjgjM9m9vzCQO3XIFMLRENr/8i/0FBB9vpMd9yCusH8YhSo28
ds9W5MJpZZKfaAUzijTPLi02WuDCsWuJScZSnFnf2rKJoMAgRNy6SdBn8lVBIgDU
3XuILqiIsm8JN6/0eP8W7DjUQgM9BC9coxknZzsrCaxZbyp8NmmmY3fZQ4rNCFLv
P9ww4Ic//CsK7+3a8IL4QNBvCl0KZ4MFb+7j/sViXE0vqeYQWl1raUxHy+X23L8o
WfxJZuD0udhxzYhFzmqrzzvg8pC56oIEbcBEYSNO4rhtx0mv6AZz23QcoB01Lg5T
qvUNoNZ6VVcjVYcl23ZC3Qv3+KgivFXikZ7c60hHPAjUfznJ3aV8R8MqHWaW1LZw
Y4RquJeuJwG4x2Au04MTIn7La9cUU/ex9KDJQVOattJYK7n9M6CXFS/z86Crpn/C
EktkfZ+1NVRtmZsJ1QxnhD7JMTvRPwZ/XeT4kiFHodst5wTtSLDKDA3osNuYJfk4
99vBWZtBLY5KxNfvi6I3t/vahm4kPZnH1BUm7/NfmVe3B+AOTBugAzWKwkCThmVz
JQbWPPl9GJ5MCEc3P+R/8EaBiRMLfAq1rDFDJZiADq+wb3+i5mfKgdGXN3RfRA+U
my87yreDFdeeJ2sKUJcUY0Yo8pAHBjveThrsKP/ZTHZ/J3wbnWskygJ0T+Kd7258
ijyywiM5dHnLyiYXYuj8Rp51EFhvwRg8A+Rd+TdzjxJmsoUp+aWZIspresmkYCDB
o61QMTSlLYLVabIBxRGE4sAT6jC0iE3X0aYb7DawcA8NcE53x2NHB6Pumfr5sPYT
Y4XTf84mEkrMb34jV+s6wB2BTyvTWc0nWMg4MpXYTr9vxLaAQpJvyHkR9tidqe8n
FvPkW/PXKF8OnXXfGB3qjnDtm6uGPvqaqpw2yJ/YLCTt1EkwSEVWtzuZDGv0Tuj7
+eleFym9UaBaSKzGCUMWspTlWCeLOlfMvgvVJ4AYWG4Q9pfMNDDWjmRM/i0HvkBd
XqQllrLFzutuFOYGG4HxeFMNrbhsBdSSw5bVh2bOgTCZY/xeydb0JHbey53giwnM
UtZzs6AVuUMguBUPOglTgHeWm00YiC9aZZm5tfZjgPsBGhFm+9Im0Epu+A7KytLX
+MANAFuWZLwAwP0BcxgLyd/e1vpM9qsq233t2S6LXGEoqwvgu9YWT3jACcnAqyoY
YMGUXBZRGv4FFTSMhQl/jWOo/e/WIIa7H5Zf3Z4JUUIG4nA+UooThnXs4I2F+lv1
LtuTgVh4gka3ln3xBpjgjlpp6vjQAdraccA9Xxc9fbsXJT+admsdhqO0411HEKlT
67sGeB5yomK6v10I24lBHUGVXRGpsVU1eb28Yw0IGB5R7F5BQF4GJyUSaA0GoBob
nz9apX8CRsLxxMk70gmAFaUI2M2bdb8t1/JuLoX4e+EExfZHbvOpa3tEsgRWVw4W
lEEcCxIyojjZPiOvOjYdWDbLr539LcI8hc4V4Mmv2nYK9y4LAoySbP4R4VfukhvD
2M32lV6fIaQ3nTqEYGwohiYxrH4bwJDiKzyiy5sF6nJfJf6sItiOcCanTbkvdI3Y
TCC+KJwXYt71iwWC++EHLLCHhDNFjKfb2MLIjaJ4SfxmCoB03fvrzrN/OcrqV9gS
mbVJiZElGFn5iXH3TFMxh+v8dKY83lujdFrPT/DiscckvfVfM615aCTNwwCamIBL
GXFIlg4HDBM+XVqbImUTZmGeU2TjHbwVOMZ/F3aP5XGZK7AKvQmn73Mmk804+U6e
ToNS7D0tuBhfHWJcMP5cbRtrKSCu0dJTCes0LQam+teDMaE94nf+rP7Fi7BGMgnf
qeyNgwza40BIxDHlqtNm6LxH4vbHXugHgMZWCQGo4Z6WECi69zLioPgSIEmWu3HX
ujc/4HXzApffn627fu7ZFI136EAOZeMM0aO9dZ6yCPV5PEoqOTk619y5AFXsI7XR
RL/1SIKJLN5vrewY9YR94JljvfGHXCRuYz3wbcmEHST6Sj9NS0Wi3VYVfztwXPiU
QujyVJf6tNXl+3DtFUhjo5Ec2xr7zK4CwLNZY9Tf6equo/ooLQRs3qpMllDombCQ
NBECrm5v7bv6w6U90ioRFf235GEIpVPUE9v/gZ8MnNndFn3lWwiPT1HGHNOZNhJY
FWRwXaZzOk/GGHy0yJ4jCljmQEGcVj3iKmIpz0/jPz30LAbyH/Khn7QogJynzFNg
5E8i70fU6daLbAhPVOaVsuQ7W4HIQHtIpQTC/QohV+FOI2LbkDXRo9z5Ev+tcy7s
VfXyWrn4aRfBA+9exVOPlbmGWR+O3c4BGVnvC+npZVPrm3UzZPlN/VFZcp537yZS
gif8xkSEMGHVRNlRdH8QD+7MiDVvp+tTTTSLy9caQDk1oA5T5pIqQ4ZqTHx3EGQZ
/atCNaAyarxop+Lcb2mtheq2sNyU9jJ7ezE4eijKy8rZWjG/HE+cn8nmwbU+ZfLC
Po5h0LzVn3zK7WfLX5EvwLxq+D+EklT3vwDHJJQt/y530oOyx6QNX/kwArhZ4XQe
iLn6AHmKoUwVOq/f9qRPx2iZ8YzNJvF9Sy7FIW8MjxuolQbIJWp4PhOlwn1zYE/U
j2TE8pV9j+8pBlQ09pPMlZzVJ5u2zU4nGf1WsrVjDDFgiC6+EwV8HJr7mpl6DCKr
wJnHoyMbxqkcNc78hu48HRdeb4QFPaCsO4s+OK0PrxWKXJ0bc5EyRzuLmg5NT0/g
XCimvH0mhocF3lU0Ub2egt/GQ+IqRhcg/fuSgBIKlNTVh4VkQp4faUvbi3C5mnzm
r+FoFjLZqDaF2VfnokGHffVLyFbz+WH0v8pA3cnezlYpSrwPiu9SouVk3STBHRcU
YAhBHBGqAC2zfvEaAFF4yXRKpaC0HjJ5fMObC/sJkbu/R92kLyuLZckCR/kbGSjF
AvL/HdQQyUuDKgvMoR2/+ytCV6LDhRHiuZDeEAIC9XR5NF0NWU8FPrfeLhPI7ZkC
0jOeuucmERMg/+7IgCngH4JdEjlb0R+ZytB3rb5WXRjcZRRPRTpbMg6CremFbkAO
zH7/bDwYOWcPc9aQ8GlK929sQ1f9gDlniXyNTFu5484cvHGkPaJxlOd4LHea1wzM
Zcn/XgNBkHCtiH6Btu6jJX7jONZW496MEGmyL0VI1BHHAlGKxytjXnJ0mQp90l3m
3WmxCHIVAeUUDw0wC2q4od2btkmT4n3BS7HfD34caEZ7EuXPTn1DraK3nDe2iMpS
cVllFl/tokZC19GVhF4368apjanZ986qOK0lwQFvr6hjHDbSPrHf9e1B6Uj9VS7f
yKTsq0aF64T7PS0cAz28x2XHIQwM/phqIursGIHmtcBPcTnEI3kAhVL5NMF/ND+j
/hroVsZRWA+OOhW5mdhM57Xnelyk6GX1N4WjXV2FPJC2XUlkO4MLj1oIKuZwYzna
iPFZw54kh5vxMl0OevakX2St1tX2qiXdHbpXXTlvKtdgy/Fh77B5fzKkeAKqiA3g
CZFlwQSQ3tzRtfescAp/7WlrfgA5a9ZcE57avn1duPAoT98AV5JWrD/0gyqcMxyE
XGv5dXnhemXbroko2r5lu3wUo2bvebNHCnLJxkdYeLckaAg/xx82e3og7uTGjNfH
keHPypr/05Do92caOtImcjUbcuaLKfU//t1nchIMR+nRBwzmfMEMYtjcf3FdpkeO
4/FePp95+Jj2hxM4waEe5m9HdG6A0sH/Hvs9EUxrcJoq7acwHRD4LOvmWNGwFcVF
08kPFaJ8q8aJ/MZpzN206Lhj9mekrOUAF4AbbShMsA0H71may9YWUwH0tXXn6NMY
Gxxt34MjAw1wdKHHyJpXRT6umB2VXbkDNm7lrhsa66TVyEvRzWbYAwpvp978VjgX
tNW5zdz4I6or91j47extFTFuIwNknCWtLKufB3krEK62LeTi7WyIbMihV62nND82
T7cjxQGLJ7ohk+VqymmSXXNbRvsjllWF4nvZRwfPvnqMSBPk+07KxfpI3yLDTX7o
0w4FHkkgwmV6bpnml6aIk1zRmU6MwIfU4Wka3XB8mEqzP4icfOakRRQ+8eN6aOV7
/VXYC3sAmI0m7FTFPIAjQAQhNPzjRBnF99XTrKl8KcwAQhVNPdMn5pcObg/RxjxV
25NCQHBpHKyhJ9Q+JYq0otBpQzDhAyB18hB14OREEn1E72hexBb1PFLOx8GAmoFq
yBFeb50Croo5mDXyPQw/va/sJL9XZJMgNsoKNVbKhwSSsxky+enqNdtcLVS4M5CO
LHJqjUBGmaPAMBLntzhhxoRuggSA8BeINV0KIRF6KgzfN7r/0BhWORrJPBGIDkzC
FC4cOrMwpGVvimAlsf7TCAe5q50aZWQPJ0cves/O3lFn+y0caFKwFIodxh+r4tXt
HVRWjANtfkxH5V1D+D4Yhxt89PpFpQLj1sFLjp9q3kQa0qjb6nKtGA0H/XvjNCF0
HuksuYbUxzcx4X0BKEjfGwTjYtJTu1Zvb7uko92uqxuWw481ZEOw1mHGPcreLWol
QAxSqJPbO3JuzxPzNNYTnxSIyctKqBzEf8TTB1H4NkB652iXyiW9CGhWDsGHOOht
K4WmVd2+r98fC5gzsaQE0xrDlwVgghHuKnTzq6jWPtJRU9eI/Nn7gGFg+ZIlthKw
9LmZhEydaJudDk6F4OdsGJV1WRBlNGWMWEuFMKSQSjudx7GFkAqg4xpPdaPiKHc5
fqvxgUIvTql8PSpkBKsSa3X9jjbV8YXcJpcwWuvlBY7rqHNLzz/DK9ZVioyFHH+x
nwja3C/L4boW58EyfFKIgLWn+cazoZjlWgJry5gTjOOD+KISlhcEgyiBJ3whA9yW
T0MQvCsVySUhgoi+Z0OToidiLuYKAy6Sv3TxR2+/kjBU6nckit6jleozudpTXU0d
dkr0o/BvVXS1eMwL8TFWzv8gUEBV2qE4GCDQLUK8zdBivoXO1HoU0mfHpDweZ+RF
zHc81Lmv/IoUyY0ShurBp1EAa/nLFfBOGrZmJ+fuZ6WqbldnZRwUMJCmjvbDvUCz
t67hfW6zfppEHsOl7uBgL7bdU5PyfPkMQTgRvPaJ6FWwcs/bgu5qQTOIu9VIpu+H
bcidGmpGZwcHaL5YObYAukiRtXF5CyUdVwkHA1+f7rtqw+d7EdNL0juq02kDUwy/
CoHQgGgi2CO0SPeYjtwI0G2kMzgaVoU+zg6GQNgJQ67sqe3WCi3sXzyItQly5tTx
W+tUEmZPP/4kLM+RAliI4g0Z3Ehn4jJqRytRYql5NWDdbgrLd51ue3IHznz04vlv
KvYcj5GRF30lHTgnx3MeWolhCgMOhirbygd9We82xaKt2/SVEMih2Q4NzJLzv4eH
N9u8mczgzMCAqm5JmpIOsNT54iTUPaAvldF4qUCWNg+CDrNlShb6FvOOEQgnKpoZ
zM2YjHxSpvmc1N2GkJM9AZQf6Yec7K9Eo5SU0aKGfRxfkCP1zVmiE7/jaVejJY12
ifU9Sytw2Qx6pbYpIdnuHl/r6HjK1YipklCTXV+PBgPJKalA4EXfeR+hRCd9OyNZ
5TGAJJCddxCgHxHxw0qo52uDXxfIDpRkiXgjhTQRFqdw1HVECv6ZkNO/SvkWludS
xX65ZR36VJvbpXPIjrjBe06OEv2uj6uPpmwd2Hm6jz0zBR/52brcyMfrjKFDb7xZ
V75aOsZE9uZmULrNU0NmJ+JvKkpsOB2dOZa0ygU2crUInCJHXvNQXKsXs6/V2SOh
yJfRP2G2OX1MIP18rdlB9aL8MsLSO7++uRZDIRSfkxCKZt4jVWf5aJFjAiyvH66H
we9eW3lwROGOK9GZHxYLMGe0g6xIPVyW5twbZLMD5YxPnoFtVZtRuizvsKCWdijj
nAT1vWX0XKczCiEe+hiql7lwfiThZ+m0K7OIACRBvuQTegN/9dFmQJuvYa1Wkdu5
nP8DhG5vDabini0bn9L70QnWW/RyXNVtKrbiOQdF/TpaUnnukeOZFtft9NNYoqsX
xPXTHXtSYO+hP94J3y1I95nPiTjqphY0SlFB+ezenK42Zxwsm+oWXxY/sjBBRjHK
0u2V5uZnityex9HbfuM3pm83kAoB+xR7BOD+lN//MJvcJ5ea8S7ee+BIIHdvCV3U
t20HNKep2ZVsQrbsklCAYI2GmUs0yIM6NBJzuI+16IR7BRihftdsUMZ3sO48LVJM
tvCrh2yy4Tb/LJha3LGBLYKzo7WBsCQU+VqGMDMvZALmh28+VUlg6oJjUDWuuTXG
1CAw3DMA1zbOO2H65W0iyiNfR9RDjgMIkwIcCDqkQnRNNypD0BAz0ImMfxTOMfm9
Gd8VYuaP4LHcvlEItkOrozdyKNbGeU4eIrMaYu1/HoJwG3HkN7F3/Wm/RnAvyxs0
aeVVZwjqHwa5WnMb04LVnYDU+JRqgT3q/V5lL7HHzCg7CNNRRSUn824Rzp9bbj2o
ItFHZIi8riNKZScVrKW/PPqA6Vwe+7msPUX5hFPrtCzb4xp3tOMaYj1hWoOuZecO
P3s+0uJ6a0HshyMbHPqD76Nkekz+BPTzpVavkF5qj58C+LDnzwkYOEGxehXNpTVJ
1PDXKKqt5R7HUKE1/E5H7Qxtl/OrPBMF7YsjgBPVXIcoWFHkUKfujbTbRTTpfz3t
jh99ePoJwxDL4UUEom/75MLCnReSst6vLnKJBDEsTYgxgpVnv1H51VzByEift4CD
4RFQ3AK1zGqPyEtJHU3lfHxVYjFIFENPjWTymMHAIhGilOtp8zQuv+pvuMJH15vo
gJzxSph9F8ZnVBktE0R8GQd02pDOf6//EuPE7mqIplPDhvyvIc35l1HmH7QQWJ20
H8Rpwo6Bknl94Bd4rb2/gD6t02UtAKbl0nFG9jsaf8wYYfXYsDKVlZq9MDyv62fX
ZaBEAEJlbBkUGN6KuZo8FEE5mCxAjrLRinh/u6h4ivi+xSRdID38v2eWQcOOEIBw
MdwkMbZD/49vRK/C5GlHvWc5W7AQhAE99SD25HUVav42qouFdbdCM5UKVSWaqaVo
YH0v1gCSbm4mZacjZKm/bSwDZDXR0AxS5m3JCdXwnq40yuacknRCp27j4ko7KfKn
7SyhjnETMo2DUltefLEIN5CsCmUiMWbQ417pIkWw3zS9IFVeyQCaqjDwPxShiUsK
2kLl2bPMORULGTX8vWgUv1D5iN+haxgwuVmF+oapTTMHb49+OWWwkwApBgY90CYk
0WW0hdVsZF763/lDlZMhPyAoaRNO2Fwn3QyxDs/V91gcLnKnjxk2p33WZ1GnLZsK
PZA79Xy260Gs0tD3vhqmZWS4uccxNFVp9jjWZ9lKuUzJHt19hqxwyJQy+bWH9aFA
7lfO6Wzo+IoT6IaH8tN71KwhPVDTHhGBkul22hObSB4S+JWIZDFZdv+w0yj0Tr7O
6EWsTRoYvF1cW6q2MSq0CsV0iw4RsHRNF8FyEn08+BJ6odqQzl3YrjC8PZElvmuR
T3gNsNc/h5maU4vM6Gdczm+RZCOyNj9UWjPKBHIVULUwsvOKPPyquT3Ops2yB9EU
yeRhGvSqwrHiEoeazh1lrHKv+OoiRV4ypv/ZrFignLAxDltznXs3kVPKIzrVfa1y
Sw9Wda2bwMjT8BQc69o9O5/3IH1YwrG7EGJ63c+ua/sssIh3P7+aSDVX8XUFbwOL
qJFc9Ku1oFB4nZtC3kUYET1JBtCsmDXTjzZa3NwTnGpL4pTadGlTDe7hmVuy0UFL
xcu8k/pR4BWLlO5lvEXriq1U5sSVlrV5ZNkznu2bGxKqadc/hyKsOw59IgoVDvU4
lEcJmv99gJK958WotDIfjLuCwBtz3uEJNC9VNwladA4DtyCwQTXpR71DnCpYy6sX
ka5wMSxFbzbIlWXqzJBbSeecqjWWvdKUjBrEPzzkbXNpwVSMFnH/pKV+AhxZkF2b
iRXjgEitRNtf6OuQCY9s8C/wOlR+0LS8IFtmiiI3ObeqimgoVdE7cDxUy7uHWBWX
tVbuaE6AqdiFvA0Cb8YyhxFSiXiQA647dxRP+hHKPsrbLDkh354YWwGj42tiGdaI
MU1zy2SZNkBX3xecS6VqhNUebk1rG3L/HWFOyFTV6SCu1z2ju9IT5S/mZ8pFIxBx
5WNocemMzZe+AFHZOC4/jZpzu6R1+DPL/5jG1Tb5bw/iUrcLdksyAlnO1nNx1NGN
XleJ9BSLCoOdoVDAsEe9uTdxLi4XApmGoGxTVB1TPVivj/NcgBIdlg6wch7ywNYX
UgusnFez8Rbgputvhqcd/koZmh9Mx/c9Qub+Ekik35+DC4PN10kuvt9s4AW9sRic
jUtl/r3GD5HDDAPIbCMJaqHQDvSq5iwKd05LOCZkTmr3a7VDWRjHholBhzVAv0p3
T4OnT3+86TeBUnfy7ITsBCPbUiBPNUab5V75NK3wida2/HmbK4CFlpvq9IQrD1Nl
TnAXYoOPvc5oGsCrjpN6+glSD7LTmNvtWJNsavgFalKpTg7LDX+C3DWUgZuVW+Xa
JHQq/uAXJ2KUaKKcPGGG9AOAE7NBXuWhqPytNyrseSKJEgIb91lLCsXNquzH4o7g
qfp/kniHNChSOKCdStTnTX/5lNn26gwR+ZmKNjeKZGlr4f+dkSRgUwPPu3jDh+Qe
ftNS+TimtQArKuhRR2EPXHoIAQ62nG9SdxNPPIasZUgaB0ThTgEWSynL5rnoG3EX
ugj9AxWpvSCNpdrtghC5YtGFb9fLzERc22eIy/3LgmyX93QLmDfDph0banfwoilT
5dD9W9DonpU2VBTxzhWqp7DKOPiA1HM4nTRhMeeCT7Bdn1x/2ZeHlgzQfQlyM9vo
2x7Gvou9rWh8XjCLewbeUEpcg7Wcc1W8NYFsC4MqSF+u3wzlIVGjaDjvy0XoZP1F
UAWI4hvlCbUivkmFeVm0KETdp4a7JYg+l53gFsdGcBaaLlxD1ty/uKYwpnEUtI9t
9YsSpkeWHaJTWSG4VZpk/3J7x34XDHK3KRCsJt6McJX+Ig2SHgFm56QFcio0n42k
p3GAzRekzenUweYelHaSvWvsPFe96lpn16WoX0Ppc4uqxAwWZLrhDJPEtKgxCS9U
aXcOj7DevHOEDshp4eAnSm882O470BzpclicRdj6Xw5GzsuyxZVY5WVno9qqG/Sl
kRKDu2OqrtYDwzrWb3pt01uSHZWLt3S1nsHrUCpVl1ZtlyiFTdk+JusxCsW5YPL9
xJpyDwX5jRReAJ+fe43g0eSaOuBoUiLIOTlKTByvmrhUW0RAM8B3VW2W7yLP40C5
UQ236AG5+KWknNgkl+2TBh8cME9vjqff4xLcOldHuhkIs8rGXqaU0u9lvb1/I1bX
jlJTHdGroioUBjG7kXbTqEJLO7HyqVc5O2U5OIioAfUYWt2teuxstEN867xFRGeZ
2OG37MpNdGCwBEVPBBrbpm4nBE0gF7T5HLLLeKr+EVf53UotNTpmzBY4e+Pa8iSa
QdL45+Y4pSVjSUy0GkYQTEnT8vxQrWlGpagmEvMHpKz7m+hjFiUokT1N6UK8Zcxc
bHJpH8bTa1Y+q1WNC7Iz1i6LQ6ZF/wYomFu9DJlsz9o5So2gWpF+6CvVdBAQ3WFo
8vQbR3tQzKSlehGIWjvjV8cIJ/I1B+yIVBp4FARHv2j1gdrAn4WC6WpnLeknvJ5c
S3ANngzVqUrubnqj1kWXQN1OpGwqbUE2LQcdQnEo03k1PIUh56Urm0az6udIm0a3
JSAj0HZk7tpfCuVsRVGRVaN1CB8tsO4epp73NH8bNc8q/iVJ+tvVTcn3/zk+gFmG
ZVJ0Xl3XetAmKR5dJZv8R+0vRnTmU/eeShtcD4EoSKUQRYUTUd0dc+Ns+Hq5ml6V
oexJr2h54beA6nvVwe88cd7/K7aZXzoSI2WRxgpPCGxMrECvtqgW5V3G7opVmAYw
uVykcb+Tp850ISTQGyfgfwdlLDhqmxoLO7P9SSWyDoCLMfz3nYkPiK3+ByiwDrMV
gYmgkDg1ADKjdGarSK0JDLP0JxznI/ZqbxPagy7HrgCEGr570nUQ/F1GtoLN/mV5
+7j+WgChzFVu37LZCO9nWsEcr/g/6T2I+WWO32LOTvnKCEaAZgz7eJNBfpP6Ysdr
I1jSSBVUypAFvtF6JBIz9PRC9SMQSKRSsoOvIqtKPNRNUAXTwJHHbW4FvcXNwRZV
7ST2eIJS80iIJ0gz1MTCLi/DW6Y81D6pTXUZzicGQOR/rfY5Nokwy0ZfxT/F+W6R
ttH8xpwfZwBoa63A77WU1vVc8TPLb5Uc+0XW+QaVtrP3yMulbCiXALiA+ofw70ym
YJHI3dC0aXdZ11e4mHTw4CFjg28xWqEIlx+xs4hXVJkGjSTheZ+Gz0JdpaMqIrUH
/D6At7L4Ks3QDyB5N2z6/18adNVxd0swvJvZBErFMnnBJVkKnVrRnrMTRUy77zqS
5gGT07s5BYFBK5cuwrC4IjSLcMgl5H1s2fBP21tefTJCUCs4/GGxAXRhXe+yNZu9
QhynbCp1N5T4MjGph/wLdo07ObTybcMbSGoLre4adMmHG4OPYeHngeZXwKKc4diS
Xzlk1tUzi7AdfSxN6mdySvWtKAULD0ncrNbB9974G2DNH4G1s7HFB4oZ7sr40HF7
L2hKlPjBKl2EDmeSg7mJVhBkJToNdPqVrGgqYQfqRKd+ytFRdCEXXiUJReus7tbi
yyIL3Vch/kP+KLZLFXGmkDHAkU3lAm3g2QWVMUpY7ed/2Nq8QmotPR0TIayclNME
yqAg4j+sSuy14yYDH2bSB36Lbp6SbcSnB/47t8ChrZoxQENKsu3retTF9CH7HDNk
BeHBmUMqMF1iDBYoo1pjDtRgwCU8aLSIUYdY0RQy98bLHQ7iwSIMJMX42u2nSDUT
MckaINI3DpbSjGSVn0HDc52XXl8h0JqmX6584+mxAuZTR9XFuFi5WYmKaj3xcqwj
Z4zxWp2KcpfysHfpzmicZ5BitUr2VSbv2QFe1O4qJxG4e5VUzUTz0piNZhY2Gsoh
padMhi5YRSVNDB0vIqgKexlXy+/17czBoqFqiflE4zEm0qY/f99MaphEp42N/lbt
sBlByAsUDnS/6u9tScNp34KHkykWY+e7Ep6koTVs3ezWVDXGywZt2GWf25kmv1qb
m8K3rbbxytGH+jN75zNaqBdunXUFUVVUCrijKQBif1X2asurFu3YHpE9qoQgnZvH
9IfyyE4m7Xwo9tnsjRipfeBzE4q1VEBHl3ugn9UAJB5epvtWbIKuBES2dtMRsyPP
AmdpTP1Knx1NoogrUg9J2zaaVOigIrY+NzdbYK5uYR2C/6eDJaTGz6Mgc/+bAGpF
HXePzUYzpfsr1uGg0Dr3yKXeDyLf+G9JXuAwEbweCheKbVzdO6IeSLoSj6FwGJVI
QZrtQZ9bkZJVJOC92fflmPAlKBGhy2acZEKPV2tKXfeG2ySyU3iB3n7fnnSY0iUn
Rl2tJTWUgGQBMU7zYfTwmHB6peLjIc8bEkYcGuT4zoVGUrtiAvA9JJx4Ci95gebX
ahLSXthOugTOxj/epqTOBg73rijBhXvOr6Ci31d1HDg5PBLIhmvIbCdgF0wDb0Ru
51QpdnrtdNPG4iPXL14lMeuAHXokeYatt3CWA00rdzkRGF4eH+zwp5DkMAJYPgoe
Ck4dDiwfduVqcRmZHyLKHqo9L80tOaBZzJr32p5AbDYp6gzP8tmNYIzuWihc3Aqc
hi86hNMZNDkrvmKRuSUwKFX+9oNm3z+Hd9J+o5p0WPanNwZGpwSDhoPoDsfb0KRv
6B4lClG+G4kzAUiK98GdlYPMEJyqJwA+o9tpfrfINN3tb4Q7gA5CxPfZLVVDZ+8s
yF2qSBhBqf8P3tfYoxRC1WH7Xb5uNbylo34Qni04XKJAlOXbDOzlGFX52W0uhEyy
D66rqRhbHaMiVkXFIFrjm7GkYTUknPUqXbgA5VohbWQ2o5UiDjN1XByWVWIBcRz5
RWgqkwhU2WVPrxxNAjd3a6zObB+8xbt4pJRnxc1XJeDG1iNx7Wp/sg0NCzXTI8E1
TRZII1LrUQazeITSkwlMcVReObHzuN1phvp8G0lqiHjWerJFoZaidRuU8FSEmxYJ
xCbqWxFkH7gfaSJnF6Jf986jWXNGrtw2ffUEr8FuatEV9e9QaNkUM4REwxTILki3
bsK1XT757Vqh6bnLrJcJeFEVmHBTWkKrA9oTFsZR35O8EHrfAicg+sj652lkmhBx
OfYqQR1f2s6+n04iMEAeyMKf80V9xftTMUkPyil2PFIAB18cZ49f7bSHqqliVlW3
u/gt0/zikvNK4ls1j7NXWj7nlfYp0CvB0nbz36lkNmPGNj//bgxVe7Htcqr3xN+r
OTro0cDMRNe1oiWdoLL92Ok0JGqzG9NfFFocIEVomuNcDf5Fjbwo8Ox8DgCSf+M5
Ua7wR60DCM3xtlVxNq7ZlDbs9lkQMqc6f154XiqrgVKYVbjWe+IveS196KLMOHcV
mLkLlBN3LTHIkta8HIOc/8DBclwCJZfsfmzk9MLS79WAUk0NVL/NZMNuuK44emCC
vd0pL5p5l1pUQ3J6IRMP+Y50KlFKsCgA01qqvbwKzQfkvTuaP8jwdPBn0E+4dllv
uyfTMyThgGb32t8SAoyIJGBT/Oe63/jpkHN2Xwq4zBfVTt3q2hdTumMJP809ruvA
3ebLURU8qOZGuxHIExZcx4fbR5q62kA3U3ofB35ED4rddh8sl4I3xOMNgC5rUsTO
/HmVtuQIySGuRYzug5BpWb5tcQxcZOaO49LWrsA6Z9qux1AKGw/zcawEA2qEtdgV
7VuzrOKfpzS6iDwl00A3/TBgXUEhAt8LCybaT9p4oRI6yNtOKwJVJUcrwhvREvB1
+tx1OvNeLH4rw+qE+eNnKi8NCJuLrvZs5zZFfEVPVpp8b34CIUZveh7vcSigGhjU
TYiGnZn2KG4sb79L+H4XSRWTg0R8qgI/JaMyly9y7LG7Mh9LU5ZJ98LklVC7E6hr
W1NMQ0AdPGlFw453AqnPqxui+ZjCVvbBdJxNGSTgZWfgfG0piJV6Jz5oLrJbCcmr
z1QLyVXaf1Ij9wCjt5eF200ymuZVQ5Z9oalB02/Rvk/3sS5GnRj91jfxcetkwuLR
zz4YNfBr13/WovHV+kjB/J69xEcAiYnH9rbPrldGdz+iYQ7VQ/C3AHPIrRBz+2aJ
+/lQkWf7JcGyCW4uL5RPvV+yIA8NYwx/CEuzGahWVwpOnYW1m7Y7yZQJBG7D5Cfe
0xVcHCgtwibw3Td1hkFM71Aqx7WW5D93zMC7ZO0Fm6t+gtaMM597zWUFxpn2zUP6
JkvLncSpP+97nPZGoGiLms4DCt35LpcOJANRN2YPZWTAzlRoGlOIyJkYWQsGpSaa
fo0CrQ0Ll4a+tUW6J+6X/mhWVL8DTcc2keitywChVr2OfaEayTEP2zi/ffrrcVHO
3sn3FY+JwwRYKGwJxYOEpYuDYdtYRfRK9VO04OXAsjyA4Ywgwdf2UboCE+pnZADw
AePfvprkbMbiEShu1gMJAOUrmnB+2bAYiKmA+SxW0R73xO5c8250Gq0NZAATRW/a
Fgq0NXF4eO1F3w9ZHLgyCG9Iqy+pccA3w1MjKZTQZhrqGva8OuLALQ9NN8EnK/yJ
1/P1RZHX9zpIYGlYol2kjBjG9NYyHWdR3YAIsUMel70T1EnProniwSl8q9g+i4oo
Um1lMcjNX7H7Gfu085E7cYxzPs3Q6HF8lLEmtBTsk3U5HQ6MUgT2W5or+VPcqZJb
uf3Kg8vxuiELH4y+kme8wxwYOp4xrdYubDDzOxYSvfV4UCPvDtKrpxMhGGjIRpKW
gUbbjdN9CPHxQ2IRKYoS3xt6BmskzO4OLfr/f2NTfz4CkC7NJFF8dTQyrRpPU0PW
oTo39UXCIaIe8AEaCmH1tFO+znGFGbgF2A/SfLat+qHmdi+bA644+hi4BtGmUNwX
HgKNeiQ+Gq+5gZBYsPS0oW5Iau5g7VPS0l+j4DgzO2dpnI8LNJpa7I8J6h7oEHEI
SX/sG88uVA+Da0y2jezMgrxJHouX+9++z6r7f9ngrfTuJLgt+IRAE0MEDXd/kAzB
o1KV9/Pnl1u4EtDJhSd5P+mp/xmhN8nJ6jl23ey7SaEctVX0nLimnIBNmShgOBXm
btacDmm+FDVW726aLYkgCPKS6S29dLArPUYfV8/1i5a4EUXKHCtW4XESJPTzvgx2
AVEQyeipjyMRPlkEarhEv7PSCPi0hfZ5ClWWa79jlyHVz5fdaDa3kYAF8MFv2EtR
JyRWg4T2qbZYoktuZ53ICMgbomNHKYG4PgcP3nVN5rFhFZpyALzCzFSdtHqH0aj+
l03xHbOUiPt/2qk6iHJH+drvmVCRtcFZNHyy2sEbRUMqr98gyIKS8SUoVWpq5V5x
XBJRKxWb7aeVg03qI3Cbq/9FoVCZPe8uqoaKvNeRVN/23yo10Zi3ZLAeaS4Mlgyt
CjaLfMQYAWPf6IyHaZao8Euf39qCqy+rbcVlDU7w97dm3C6cYWJW9HCfDEZbMcWR
/C3QUbaur8p9QX5UKfeKnMeFRONlLtEPmIy9m+iiM7MpJGAo5ksjO1BsPQICY3bu
d3S6/1WVQdpG26aitJUGvqHuLCMxgrcjY0PS/uiG074F2AY2bapXEis6jURIZWuS
36srQ38qlSFBAYR5ltJl1CaBdLeBIy4IWPUx8HhRKWm9GnQJGzu4rwBvwwGzdoL3
erWBFTF09Xo7pzlUya7YlE5mfaw/vyMjJODfC8gYhNoImaFYEyH6J4e4IahDM3v6
B/yo5sO9fRqIFo/E/ORDNPNfrqT5D62ie3ukva7pWiuL4F+KqPKCIGfUnZcYzItx
6bfXGASwI5AycGtCH0pJb1+wW7OdnyfA4jcOwGDlVrrbpC3jjeM0aQIdKLN6bf3l
NVhoQFfwIt7qgEyyhW+xs28Z5oPl6QCiL4/ViqTZnRRwKUBNWxXfsUwghAJ4MR2l
xHCJXeAQ1sALLXtUVqeiIzcG5kYdu/4tLIWhNNLxNYJjFOq60bTnbZcN/SD7Tmz6
yFw8q3roAVQ7S6faqzTewd6pwAqS3gWenT994E5MtpczNAF49GPAdz8eMMs3N+Wn
9BzwxT1wjQ/yfWgaZzbuc2DhwRkIHbxLFSpgBU6qZXkhl7qSNFB56zsYvqOSGQrS
TE9EsesDu1YoMY1xDu2vfYdnXrvPvRAZOflmvPuK9ck4It7CdviwJqB+Qi+29nyS
+GJMJrYAHAQGv26IZQZdOuJ9gRXTvV/Hr719p5OEwm+rrQJxpelGS1N8OIIh1ZST
gpr68RXaVtHXejwgBZRa5Dab2dRL39ImgVzKBwuBxxU5aaGnrJntL4JJlmVCZno3
ucehDNsCg56gZSKhivPH/ntCTtfshuceKRMnw6Pu1D5bFBLejynkcB+lclGvbFX1
e0mG8rxthP/y4CrSW0OOc8mM0aMj3d1fsfq5Hby3V2vhgtX9dOIcR6Xss5XP+f7v
3MZtcRYOLSmtQymJu5HD+FeA7l8o4Ty2xUosaeWPwNjasaQL6RroHhb27XwTUxrH
NQrQS70HlNtAzr1yRfY/Juzbuf3DcfjXpwuVvzjtd5iKq8I2Kd43QwzCXpMnusiD
xpLqnMte79RHzH6FleyAh7uE2Aqla2NhZRvRQQJucDD9mDYqCl91cKMMJJezWAH9
yf13nf/jsJQInqW8KMOx17Eye0crN2NuLUv+MdHS4RTlojPBByEyF2Wl1vKXGaGi
dVcreRgEba8VKQm/5e5ww+nc8VsF9kIajOCAqHM0TiRC3Mq4XVgrf4J+oT37CcLS
mLdI6J4HfSPB5EYJrC45QjI6zV/9L4gLgh3nRCvEAymGb7YnRUOlR1sI3Vh4l+Om
4RByt7VSi7C2ShZD9+/Mjy41gkWcXORMR3Z0FCjm/YU4Np2NX3SRVaRiP6GEdVuo
wR4c7hWWDRcRsE5VIBF4yX5OC+m+BKnLEFpeT/AisfXP39nsgnVln7e7B0xxCIQt
kegsTggGI8s9X9dizAppGw6Zm83BPyVH3YMB7ZyJu4EBEpwlVpin8eT8lK147g38
CivrKabackMRONUYgA+OG+o6Haigz7c2cbkBmnM9PF+dUzXhGaroI6Ky8eJq2hW3
GpaI+psGBW0mnKkohUCVbdPvhhsneeeeLUs0OA+Ohg8oMRskXddy3uwpjp+Cebp1
v6l0hu8k2ssY0r4ZP6KSW/Gv+Jqzt0kZtOwDIyT3elrx3hh/XOyZhX9VHbjphWRb
hpF74ZHFpC6U0JXmnclyAniVnCocWEdZYAFzp9TVnSk8xhz2tDX8WgU+Mfyo/nPz
dxSybrSfgm//3pGwJKZbKKZRq2YIbUEJArrzgB6gL/yFgHMN1dq2vwpnG8jVa9yd
1JxB4yVS0dWS7M4W6Bd1dMKOM3/h47DJ4pSfvjTLaWnmWbLVcz71iSFU+taAb8vt
4yKjzXQIstaX5oQvBb3PD99QSh+fupXYGCfMzJ0rarqOErk29XiQhLAtepsQFTHM
yKjX6vniaMDMyo8EMc1GGz71GO6L5k7w7Q9VHIS2JEWLQMShuDyoyG9iRDJutIuH
S6/70D6ZzDse0RuErN5nsBpHspfvzRp6yyjXOzMBoHKLAqh1631c5mxeE365g+Za
0Sl2ZiC4D9hRf/vsYHXLR91alo8qBLmXB9GpW57vwgURBKM3nHB+GGp6hURKP49S
ymmkdrSpB9i3SPcJsKVgpmPckBfXkeWaAAcdsB501+Kzx7dUbry4FS+V41Vd8tfs
nvmqscfiZtr3/+Ni0NHwsgg/g4EbZC3XuFu24rcZEthei4RFmBPHVWv66MxxHdVX
J+pDcbw9zGSDCoAgq4BermtqFoU3dg1CRbxkPtizQt0P+JqnF4bgH5+6m1PHAy3n
syd01ejEmqDoVDjb4jf/M9Z89YdzpW0Kg+wb0ppARxfHHUUa0IjQDsIP6a1+KxMb
23cS9w6LtCFm2UaOm4TX3VBsQLz+080Hs1t6sOvCz9Z6n/GRNpSR7zqOyE5cflVR
mOWkQsTdI5zOTl9mCa7Pwr5mpp7oiiuea+1cYjszCA0bf7/UBph/fWGeLiLQ1YX3
Gp6XiWWclvK7oHAfPBINpWD6MUt2dUkkKzKRu0FadVMUIIM2UGUYFbyiG4V/X6n/
5pIE/LxBDgd2LtzN7TAxWsdMKgXitIzOeEvU0cE3Ta2R1uVpnGpyQpn7KkiR402p
RZDc/okcB43aVmqB/BWwnWfjWLRbVib2woe5NO0QwTCM15b4nzK2Lxa46nYUbclj
XvH7WIwbY2zfsdIoC2DXhzfWbQTGvssD87UMTQcy1KgMsHywS+34Bb6i5CYtEtd9
gx6IeKb9+pMN3ZtChm99s/Ucco0WR4E1IHHkSCaYMY40uYBwgXMUDOroeZavPPnW
XE2uUrrrPRlNlqaGlVjL/CcS8ttPb1yfcEWFpon6kFMXfh8ghZPh3tM53e7+eoo/
yHX0rzwd8ONwXkI7g2U1mJTEpGPJvi9HOJILudrXnmdcr7q57IaGFe2B23Ykk4UJ
x5A8bfC9zifU+J4cutXkyceO+78zqv9WSnmu24BmsXy4k3kbjqBUmf9iIuv5VIy4
OL3LyUa59mq6QK9VspwsP1IKgGoFgDvjPZGO3PFyBIck5maMYiPnLDQLDbDHTmkt
adlzfIlPg1faPMDlLeVU+dY2YDI8I5bffB6AlL5nkilspe0D5Bkthuc+/MQ5+WyD
npRRZA5MpTqwfQE7Gg0HKmiHNuzVCi0hrYnHvksM1fs0JwFaP41FQGyHSZNVP+Gh
odXbczosbqkxIFSBu8Cf7KsyDamhdGUxXagMS+QfLKB7AGrBufzg1zhUf0DJrPZ1
Q+HlTzy8lKvNZybNzdU73Xho0LL6VS6dphj8kx0pkJcbb4jfVm69Jgkug/zZlvId
0i6BaFNR2oqrgl8K9ZX1rrTL7P+W5TNOsKsntgnmkRf79FtqXAsJ4L5REKPT9lF8
Iy/WCTD4hQR8bt/rz4reOZ5j9THIUmqc3P9DhAIKkPrzEugEMlHSbTnE8UiAcTuA
SeJyUWDlM8Jc1WSvhpUnc0cGYvxam96Z4nCm5RMmTzbpcegzBXGuJAqqv5X266ep
BVFie8fHdrylYXMOmQ4WOSU77I0ReHiDsQ/7XlgFewU/e4qkAcG3ZqHrmLeyy15H
+PVfStWXbz4Ml8J17Y3JEEOMRxf8fvFzqb83Mpr0xBTtf+kMcrpbAYQrEqdo7hbv
+pXBottyMRl9c5j5uuI7egelq4qe2XgyETNS0KRIunMcp7LQpucrYBxdW8VaqIxs
PnGaoLOq/AaVjdrUy0ZpktzIVd2PycFJpmQJHF/FtuRqt7JICp8svGHfryX6LtQo
duyuNPpE6p/To5UIn203+nA7i8nvpxRyU1bnAvqRlP1X+j5BM87VxCNwpC0Z05RF
Q6njHagV4LrqtuFB/DOF2t/Mj/8YIL5laBMQbeHOzhEQUInNVaWoRf+selyA2H7S
XjS/qSgZ48xYECZ8KzhRaM+IFxiQ1EmjfwHP95WDsluvxnTQuMXkubUOuNwdKqEw
DQBj8tyL59r04e1J2g5oIKTOOJtatOup9CaJ6kif73mjM07kYMLKgPGKDcuM6Ny/
UmU7oi3a//C0D+r7gvxLgjht4Z2iHiE+leqgR1bWC/BvwhheAr66FB7qRTuSFdeA
ICT9Weg5cKeh2X9xtgpALqJbKD0yFIWRc16I81AgXCn1D3f5rj551EKC5hBwfQef
QAD5TsgwrkHPwFFKGCN9qJJo7ZqknXs/YV9w3u1pWGgMA4nTJeFM2oWWpHeumq2Q
EuAgmG9IMY9c7Sou/cTS0jbXuwcvndnDSagf4TKTSFTmesksCM8JwJXrmCK8LA3D
GKDuP7FKqkikSmMu8U1zjtypZvBaIPQ9sXF/51AaOTFBw3fjyHKHki5b2sqGgFPp
AQZt6oW+fNhtlQGgyzi1Io401VEyOtbPlxV5pDDT8TnPiVWTWXNZYDMiUQPiuxX4
CrGIWDKm38OFgl2tsKbmTWgzwyx3lR93tjqGeIorSgOsiog3Z7yqUCFHyLJuhwg7
ZAVFfZ28estZHtnduV65pbgqLazK6U6KoEyCqEN7y6JkL/vcbbnyTxic1aFtV9uC
nMtNXsd9KYh5QwjWyfgoCVWIPIDuaZDIBWiB4XaP4Omzt5BR/POKmXwI1J4NoV31
1D6ysoGA4i3jhTEKIGXflYYhB6KHxIfkkgLaPFvcyaEgz3EOQEqAX2qdQaORxnTm
5HXpDB4obxMNG4QTd7kJppN7WpVfRTEcTCfB8ubh36rPyWB+CpfEvUmv/zexlSPp
ecB6JFy6lWHh5LuTZj/Oxn/CG8lHKdjAtFC37S6zBvbuGa82Iz4o1NXqyv9/Zxh4
l3rimmzcxHwJp1p+NEvc4Zf1JMJpiu459E9yYO0TkaDNqacOuvjqxY2Z72z0LMb+
cayXzxgqvbTcwyGVwtVHeWgxTUJ7Y6a48KUbt9bXRCIGMaS0VljDnAZCJx+sY8h+
gkd5H3vd9tNk26zbRx5FzCWTrGyoLNmzrkiKSr3iikMrRZZxxcy32pKj7Hemaqpn
kf+gwKVqUpBjgfigxmjJFGi4QfDaf4ZS1tDWfSuS9LkcQ7U1mcSJnGDT0FJuq94B
IAGOUj51EJNHFoOtt/LnJcqOgbuCPkUlbIgGhHqz2A2jhz7e4xQFpE3npgv85obu
tpyyjMHG1nGcnL9Jy1zslbbTpM+NT/ipdFH3x2VVe9LonTyH6O7VTUH83vJeP+0B
rA6SC552SmohW9KCq0dq6tHiQXNhs/nLPIZpXJSQfP6zDax7XHj9Tn7WDqvvaNe6
7I9X/S2J+svC3lFghzNf05xwDs80BzWBeW+o3hMsZIDY6DeKE79jNS0CzEkWbQpa
1QRk3LiTPcyJt5ThZNJxJe1VzzLz3q/iobyvr2QxUre7dV0ipn+/igmr58s1gOlN
4n417/ixzK2QbkegT5f9BxeIjx3ghHh15MrWVfhgE0Ux6BxPD4rbNEyVDLQv2sw9
GtlKpU11yazvVinMjGi2+w6gL9pzuu70BozuKoYxFJQIqdCX6pg64cyrTcAk+kob
QqkymW+t3wYbXutcuybw54YhZa44A3tfgzTs+bSsJYoBcFvmujFLLKByypr0w8t4
ahCJNK62JTWQzTySGwjdfXlAOZEjefaWmDFH/1MVfrSRybj0o076OjylG7MUrejx
LbQEvSdOQ+GZ9WuLQGrqgztM+kILPZVE30ADXJ6jSeJmH/5p0+1jlDbYC+2JyL9t
uhYKgR/flOdT4hS4az4HV4wQHJUqT3GWDOp5bEabUgSN8PRodMd3rfn8KM43n+ww
R9ZG6SwP0gf620GSgoesFugFDsPM7Npm+YkjnVGs8Nk0SBr8kn29Mi+aIW5WeELF
b8MPrPv8C8uYv7+hmtYaXxg8+Gs/TVq6P+7FahvRVro6x8K4IAE14ZlW4I1P8B4c
AoS5zg0+e4ThtuB9i626F6d9K1+XF+UhPA5rcq9/ypJb2SwozYLJchz4QhZ2t4Td
wl2E4DVlYPXJalJ/6IgKqia9TKTLyryt63KZi3/dCxJ99FU1WtyTPC7hTrf2HBvI
QjNOXeWq6Zs4PLfd1euuyU2C5A+b5zl7lIIgsHTik0SevOT4guKOIRsbYYBJiMjd
VxP5k+RalwSIpmkPX3LE3LPEwZVD146pAq69Xgo4fDIgGmRTqusgrNzrL68t5tyz
yq0f5sOnkB6e6C6ZXkQQs3JkaX+UTU+F08HjHKB9U6kZJwkqDuLkojgp/JkXyLLK
+peSOkDWKSW+aL+TT4JfkkTtPweV8nnkXlHF3R7LKbXf0Z4Sdqy9RCyerdDQL1JD
b7PQNRNu9EbFbhO27xAYgW9yrpIF9/mPEoQXL2ZV1k70m8LNXEESX5jvotlLgRva
wEqyJn628m0puRduuCsR4IkWdaIb5cMgmIQKmpi7Y1Q1k0510hxqn8D2b+Xnl5Zo
OZF3w6HYlaD71k71hvk8XxEP/zk/xTOHpFjBtgp5xzP4t7gjC2BmSKe4pppglw2a
rhwOTUHdU67NDcRucpuNMIUJbGGd/+JmGtyLALjDNuefG7KA+vKnPPA3+OWmhdQz
scabwOcDn+JFnzgv74qKPEOr5lYDi/30SGJvnstg/xQq68wRnmVSPLi7XVPIjKRZ
K0zDTgGO/dSnbOHi603YcteRsC1Hyvr2mItckB/tMeumTt+GD/U1sHFPPHKKdca2
Qyh/+ugxDJ8Y3UAiMfB+ww8HSEgP79SKjkhWbFqoHk459EsLP+7oFF0T71V4DqMd
2DdjYpr3mU755f9vd0KIhPqexm5hL9LjjcDmgvpbbJSnDryrsLHYI7Oyy8kvdqbz
KXzET9KHkEloU4cKWjVlTkJutErQKapi15qjn3gY/GIZ44/LhctkX6Wv7e/HS6O+
v5+AThzAFR+l9zGO4/6aGiqS7T1nGoI5iSIAne4aEB2RyGrrEIOqJOJ8Q5ii0736
ucJbRlUN24AffEZOIgRrHzJYUycYT1krYaeJlK7zYnFMWsOsHYRkCpMZNCvV16BH
yyTYRTuSUyh/YSzSynZahaCBdGoCCeHWnNg/7YFFtfZFG6Ub0xhZGCQRZt17nV6W
MExYFfLzw3B32efLpl5kSk1C88a+xvoFs8P2GgV26qBfLa9sPF61XmXFcmlRwM83
OFFuG84HVAxW6YxrFTB39OUuZgQq5Wn8OaQ9CQnEA6Q54wVqis+YqG7irvmC5DXG
EbOBiKerugcPuEt63cI2K1L6l7A1gpXph9e4MI19m1Jy17ul+yc3K2mMSxk+3/rL
SwIzmWI6M5TqqYpCZpNC4W9wWz6uJI4bYY2OZ3xzXPKq+Jhc4BUEwL03kVRLv8XG
UXEHpy7EzhDdTn7TXnWC+K/7sxujpzU+gzChhjBwMdTPq4ova1BzDQuE7Z3vAW0p
FLuTKaSYValP3uvpQ1VClfJ5Vx4lzGGKpyCUNck5wKK9qYIVnGV/3HYixUvEKdND
OzJkmb5a5n7pdUlFBJ1C/1U6o1TorvBfg1tVU/D636SjLUlTAp7DyP2G+3ZfqXSP
O8w8PfM7j8vAk9xT2ign+34jnudhbpoz2xl1ETE0C2IEOh9XOnQeggantdY1roGg
neR+Ei9bgSVFrjx3sFMuliZLUMcQ3+JgVV+Phh2Q/a4dl6hjR/4R1vc8gSl8KOAS
laaRP/nMyUA8tmSp3pk7y3YHHiLulgF2OvQ8/kOIVyvoDCj+IZikogM6zsuNcyhs
TFiM1Qfl5xKHywM86P21SRx0mk00b8rU0LdQLI88KZ8Iymz3WzWFTVL06qYSrJvF
BkTXRirNv4Ab4nIWcXSeW0rHmVEw1b2rIDU7A7D2mlNCFNPR7uNEDgt70ZMCQ4m0
K4tt++yDYmPw3ycyYOQQ4u3KgqxCEgkIIuluc7g8DvxclrATnrGeemqC3a4CfkGx
6jUhiHPzUKki26IGd3u+F6SOr+MVcqVw7r7JVOm0Qa6cwR3zK+JLTxcVwcewWH4f
tG5ZQve5RBtBNGRYj9sagLIo8NBhACFyvoFvpHoWA5Oiq3MAng3waZ8Wj9sRwR1l
jH4kEC/jhuArZzHuXQVRhaUibxdvxYs4zt8slgfkFz5n8Kph7w3Gw+KHV1W+sDWS
Yy5J7wYZ1JnsomQd7GnBm57nj7T/x5WbbKn2G1UvIOqwFA1rOMwWCjGD5X6b1wlu
pS4Z5FtjfAZDzsCp5Zq7r3jIA2llKzVpmIKfn5MIbe9XSxPxVZaNDqgPf/WTMyRe
97zym7FrW7neug2UOG9x4dyLzF7BS6bJGSOu55o521cSI8PEiwaf3dyIvFmaipAz
D/MgurXQBC27rfv0fNxovf3wACmK7o0Mb6db70No1otFXF3c3Ka9uddpCcG2RkpE
7S+7eFEmnAd7OyvigZjumHnWZIj4YZ4ZenzAssfRtY/5e5kngT0XgJlC64eArxwn
B1GfHqTyd/zKukTPJlDl2yLmoW018CSW2oTq0DnKwDVY4tTSIydTdUZNFyK0tuo3
s86P9mSYA8YMnmk5ekfknpCs9msJHZQZhCw6ipE0185MMv9MMYyA5UiPyI6cg9KY
8nNhclXC1PhxUfebuFIgMtxLZQcuoBafnzJ9TQLUCUCml1kJ/DTu4NSTBqHWBazn
liOBg057SEBKxAukFJnkqAG3wsGPbYBK4fcbb3hkJ6u83LLqKK50Lk1t0dDDfckX
rTEJFyvGTswzHIxnHAW20B77pm9XqWiNnc1WFpI1NG0JXTQtYItDfYnNaAG4Jkmq
hcXAQpuiMktRmhYQB7iG0o0tRjTpFFkTT8CYWAAKCdssr05BL6i8fnGYpMHwFbXo
xgURbcD9avs+azw+I+ZKOGEWd95RKnOya6VL+FstHAtgfJwLBV85Xb6ptAhFz3lC
IZkLbXK6CnegtdqiHfmarNVv76+ufFyLosjNAakcrf/3C1zcqmjW5ri3AZi5TCqz
nzuDRW6lDK/VJNWMDGb7wBzNz9f7VYK01t7Yk8iuTBlxyg/N7pjOjGi5ewf5WaoU
hwuVzolNAJ/RfDwJM3jXO2g9Y4bW5X+E7cfOtHKDydfzNwfMuHPzzU4rk7LRFlD7
kfnmCV/8e/RprvMrYYvVXRxpk5cm2AtrU8Qz1UdZXUehIDyQNjqQ+peSrSjk00Oy
KPfcZjjkWjxr/eAEo2S5DDCibgUNFfuiFCiQjclTepwN5XBRsqDViTBd/yWLUQJH
+pChrp+H8UQjJ8HfosFgjfxmezAd9yahbrZm3zCtHp5m8sQ+vBXRQhdFPvaUFwb9
Fkjuce/szfZu8DWsgapUOYuxW/ER7otZIyjxnfPqwfpefeVdcb4HPP10hp5e3xN4
qLjIZIyfPwH3mkDpK+O1oPJhmyCN4dRiwQU4uvKs2CSh/4QcutX/GL2m7LXzuecc
Tc0ZA4NmUTO1olj9JpdatB0bUEtedj/xs9MJYHSOHCJqJhwxvjVWE6AKCo9bii8M
z9pV7vI7tZEpnohsm+FdkBKJdZ9mM+eitbes8JvOZjb3cuPOQUCgOqyl97TdEI2a
100RlK2xedFiBkOYVYp70+scsIQiEeKwTDtu60DfO9ulXDFIlTTWDKQVdFXjg9MY
k3raLF9yL4azR0Xt7vEvcokPptOjuTpe2HJj4PK4ANLdl1RN4HNdEfVjammncWON
PkD8pXmC6hVrpge3XsHWAcVEIpbcDJQADJ1zg/KW0AohT671Zmieai1utLSM2IMf
1Klu+T2baG62ZlTCIoAFDPlE4xDN+IxvOtiyOQe7zr2tWF85hLUnI8CGggIr/BkQ
YPKmBWvw0utQiLlcrgLO3pcOGXVAl/eEolILLMVQfGVNDD96mCHLFRydOtcnDAvL
FfGJWtZ0IWR1GlThEwl0uRXSZqKXzlWOOxHkA7fnt8EwEr78Xb3VEUidoqgQTXsm
/82zGr3LhsWLTZXTitd1Yh0phw7Q6P4sjcVaD5h0o0bLhBiOa1wz8ImAuWxTfRKJ
9z4Cwb/1KjBEf1OKV0gqvmF+jb+EsBkas5nvM5zpryzFeKYxOf5fFn6Qg3sAZsyL
JS7m4Efp7BGSwPDh5SVsSzXXv6VxbL487fLSRI7fiJNMtRPNkOEhyGG95PUwLbwc
E73SwscwJsYeSu/OLAjHxHqE7hUT2CDei0mP6IT9nj73EFIq1uskWY7hCm0QEpjR
Y/647Bt5JQGU4yPtAfP0aU1tTRQM4uHnXXDV/rge5xkmPic4bH8HCjQDzLW2FlFU
oGWoH+7wREVvRp1z7VSn5kyam0eh+WEIpwFYLLNQA8KWxNQayQGc6Tdq9pa4do3T
ARQTLfJWa5kOcz1UujvCAM9K/2BlFtkn97LBhn93XPmAEeYNJwiiQC7S6z/LxmXH
cbhx0MtilM9UhirnAscf5Q6NsD5vnaXzoo0szZ9Ge94m15FhMULlH+fSMoQ8t40A
Fus78F9MjvulSmFhZR17JqRViIZQx9snuWpIbGddH173xUPZqRn49LgScQM3SIJS
mJurFMxpLdmiiE7NKZD2ULZZi/reH7c5fTghvyCcQJOYEZMnap4Wj6WReqSQ9AhA
g76c30fK3CuUs4Dy4PjyXWIoetk/J+JF16FmsmPUIYNTAf0392/n2AWnIJs0+Ooa
lQaEl82/cOQzBHH5tl4EdE6wvna54hSikk3MtITxW05ck4CwVmzcyToqoE3J4EnN
AOkaHB5kUbs99f1iCcg+CHmpWH23/zUjoklctqmaaOJ7jUwvrtlCAtlogmFsEV0H
Iz3eR9nqDcVMqeAh01Y65T799rFw7e0JK71AK4GsYLAL9SjS5/iuQoWi703SC6iF
gAAY1FV/7OeOkSTWUmFVD+2tFYYVRl4sk2VItzaDk1dOiQiQDj8ML8YLN4+sWClO
pcV+DOCJ5v7Qi0s6lIsDGn3xwA5LCdPW15cHQ6x9snSgtVPqrjvaXYTHdDKQ/FjX
cQS4lugt7vZtWJ1q72xBOBcRQiAuRpi1rzkLXq6yNKq+LUkMeMs5VwintzOHh+l5
6hwazj91lNfzlYFGxqhghKETUAtnBaG509DW2TZ7z7AcwcXxlnI2Jl8+4Au0Qvb/
n2WKp3x5GTrW1VBH2KrmLXJOqR+OUitXwD+S1r/66FM3exNLt2MFClINvqSNBbqQ
nzZ5YzS71e8CX5M0Oq4/SN/x84UuE/tuGiYFucAg72kYQwOZiSBWtjumI6lNiJZT
ygmO4zrKThwYnB8Ni0QWvN0eCdyEyeV5FRreWL00kg9ahnqw3mNnY/P0t3brJIEv
b1c2GmgElTaseRnZEyPx8gFW5w+EvQ19eraxCnY7gm/KnmbMjLYZMKNnLqAbwfCY
yx2SDP2o8jurxPXzn9pRyh5apQOIq4bMt6BgLp91TIoqli01M0FyfgUZWzbu9Mcd
2F7OX4OKzekXNMpD/6k1HRdtCzdyb/qDtgzfbf4NbnHLdaBeJ2okG6xESOiye+AT
ZWD6h/pGvm2h+v0Wl9D/AIHbIH/4FqLds4G072Wsbvg3p+4S8xS35tzN742AYObF
Tf2djx92Xk1XqjhtznBlFvnRMxZMPgkDz2xezVY9fPQh6KZM/ltpVUY/0//EMLZA
Yrfak5FDiID/AhBgaHJvMG9wR91SGou8CHJfokE9rifWiu4kPb5NBvkf5VeWTSci
r1D2ANGaQa4j2yBZkh4TOAQDbtsVW//wRpyCu2dN+IjpFIbTAuWrZ5mgoXKm5150
M44lWuT3yYiCqgtRAXBUIQS78wKC0RsBPGvBgRmwlzPqq7q5AUthet9ZgUhauUvh
OP94e4SKMaHxUuahDIOTTZcrP9VMpK3cU2v5MeykQIywMxfRNfJ3SjnqDxkjhT1n
1DZuf5xMKzObZbqC1AN63Wt12YowoudBxcsKHCHwErMYSQ5jIImIKjduTh/sWA87
YAXdKTuiJsmRQHpWg827dGbLKamPKODxisZjxB7/B65PyBwUIzm6PgqUEEGd/2q5
Xyw0nA/fB48c9J5Zd+XMka69Qi5KrCh1YGMDLWubSRxNx/QaXas7qPcHRJ2Ce/QN
melKeZgkIgLg5p0VcY5xKwEW79sktFDezfyxiM4EzBakzenq4+RuFtNBqJbr7Clj
X9LuTQYlJSskf3St+I84ooVDhNF/sxZ4qpzySJfBPMRNCkaf3CdKSCR3dbM4vhGM
Mk949g12K66XPY1ANDsFxUU77RnGAmLOShFGN595Y171LOef/LNW6q14Ikb6d8sT
EaVmgbtcZN+cFWFNus5jf4st0BJr06GAA4ncZ4f5c6Utzsrw6qwdaWKiVsi8p+l8
yYTCgRef9BJRUMq413fwTK8EeaAgIju3cQWGVD8QpQi3XdqhozWkgt2z/xlU3dWF
2Fgc9z1bQTGJmBLGDuJw/K1V6qoh43qBx9oLud4IcO//70UBB9rdJ3KvTPTF/bJv
ErHaU4W0dKw9HtT3JkMpJx9hmydfrwRvfwCAIkFhms9PNTPsscAD6KIEld2IlM+Y
H7fdAieBfcYLSekt9dV1E2lt0zFpKccL/QbDNDndAObtjQTe/Xs7c7pvZ0vm1FSY
eSK0AbmFTv66KLjg2yjyvr5Aoqg1XYkfScZGcm8fkPmkBzQNf4hLDPr36eL+/HUg
ajxnADhAlNWewA0K3j6DZCRWpkWg+UFttVAa8JddNK/sSVabNKSgC6B02E0kTa18
aMFXJNF0mFq3pd52OgPBnh2DoLDhLgGGeDAtWLuFl3GCs7i9bq8a2qJUHdSt42Yc
kSXYJSFFHVb8SOdLWDw78G+2vVVuHrbXIlIDxl+FgJfmzT9OLw6kGSEabGz8aqsG
IJ+8BOJ9YCOEKq5FCCxovKTf0V/JqnczE4UwTyNv0X1p+qZ3klJDjWcoKygFMrHO
4DSpHKjos1UtOpfhoAgolyg13CfteQdUJRkP42moVqiMGR93p/00Qix8bNQlIwbB
CJUORq4iXqmDiYsLIAQ3xmpL7Yv/6edZHnum4ef3m/Qk32CxLYgJyR4SrG9O7wv0
JiSfmShBspOvJhwZ1slzpTnc5DcLMamgxW/XV8TCUC9saT9Fug8G43WzbM5HnAjh
tHU3VKqmfvr46MClQGqy/hAH1Nv5gHgvx7ekmQX35Ddecg15qMbgsNZ2TGhUhJYd
8RgAgqm0z3ZBBAcDU2kESSLPN5k+SGxjv4Xz3pqsrp7HlQBXYA4dEbxfNK/d6Ffg
eVBRTNybA9OUbQ592KCkyOVHTCer6qixlIdiZFlUbXLHgKsz4C2Hy5f679ox2Zkw
KsNrUY6xEs+xXb6lbfPZOzRbtIk1rDOj+WyM6vMEQJ8px21ymcV/IvEghamBPzm0
wfjvguBFMOfx0g26/A4JHZBAyyhW23Bni06KLs705LWWUz+t6NBfNnyokAyh06VI
38vBYBCdLvF7ssyKq2fSkEaxjCKEtldaEMOWQql+vjena6RPUoZJMs8uvR9OfEip
a22mr9BcFeHbytltIDCioxlrUM/FbPAOxXe4cNFOqsGWaOA7wCrN6YRIxWLVz2Ak
dhRCWwAzYtCwZ7CXfMUHDYNOVZ+4YHXBWDN5Cw081QcFTVyVwWtIEyogeq4nk2GN
RCku2rNKFBP4XbWdQd+6wmsO/wjuOTeV1hVM4i2+JgujFGun+rhMoJbAJ6NMBAOF
6YWiihF/G221rJpDYCUpo+mHuwbFsFPaxo8N/U4JB1VNKhVG31aR/xZmR44z7dbl
wIlrFJmAboTV/NhpPmbJMWNc5AJ+32KEcxFZVDPDh1EhuebXcaiyurFk2otNRQ59
FYnujnOiqqzJTOMGtfYqQklmkR/IacBxrO7GfvrtN/D27axOuH2Tw2iSiYtnOoIx
WU4T/++lmugpKRCA7Xi7O4lyHCVjbdatAXXRBJ6BfzW/iPiET7UkSzX7C7hVKCuH
GE5ac2cRCEParDYTEjT9HV1ov+N6/S9/MfkBiHRjkjGaGMfQpK8F/fs121LamNpp
Aiq5x5A5hfsAPeof9xEBOUdOB04Xxr6cr9hfqSwt9iHodIS02d8aWaLJGjlJ9APn
WDbMhuMrzjnOvnnEl6bqSua+07AT7V97Uk/2f041tH3ZTcVekIljHyrO50B4Ql+Y
kFd6clCAKYA2QvcabX/ecfzMyWBprwZTGx0S4C7Z8YLBRGmwJPnBgA1CKW4oldYY
k7w/JGtSYeex2aKssBCloSVOGDWLfx3kOvRo94vlI7xaV3QkQ/gv5XtnESTgBFFq
V6/U87GHfIe/vSmyBjtLvCzFs+I8woSrX+i9qTc3RGtt7Q5JDgV0Xx6LymuHQKPe
0ICT2AdwLJP0KWAIJA/IxoD6ZLMDMqWTfEdqsjMj3DNFx0GWe3HgUJAZPzi9MaYp
Myugfu0LHI7BAlbO9QM7m5ZGEWHlcNfghSfZ6ZG/9aKo6Z4fgZzrUFCJmPhX5bck
D+Pe2e0ct6c75CvOlbYYPRtLTvRsleXG7bSzReqchmHbg58NM5Nq7/eTn306Y+QI
GSROg75xMvUa2He5m+TYOVVj8xbBZg47k1737lAFqcCxcj63s9ldbA/nC6hUF0Rk
fH/f9SHdkWnexncRGDSRmYSS6Jg6JpI9pkKMiaO/9j7BenAzLZ2H/tdeAxN6jsg9
uAMsVs4Dr50hsZHlLkRrLUoQPJiuAJtPdbxsfItb43DRAEY2kZfL7Oj4OHL0FhE1
JEDDh4I6QHPxAEOr8uflBLZvmyFc5667PFA26Li/cKsG2YS/2ZFcu3QZqdu7NvYE
/MqWJ09ZYJ7g5iQdzA92Vro+NIQduh9LMIHAmpgeeBWJB9vW2w7FM7sgL1bzSPu0
zTijZvmYzRvtq+rfFvZhn6DxTgvtPBh1SYQxQWFGRok91k6B0R8vQgR+QJr9WVlz
XXPFp2PDmfNhbMHan5n6bsApamS8sNU36bzfHn3aNjdbSNihEv+0ynU9ZUWP8lsf
8Y9feR2ncUm1x8YCeks1ndsxaiWv8i1kqjZmep4vnKFbvULoSKE4ansUbn43dfw/
gDCrhDKQmMa9h0xWT8KTDfT7ANV8jGFykZ7Ib5nRldv1H9Sfhx4N36JXe2gfp+mK
5YypDleoSdWxUvk6EtzjGg8NdA8kYlCuQSFEwZqN+jUnhaj018QAMvLzamLfB0HJ
saSQpBlY7uY8LcSaxoCfDfAEcnqj1W9AFi7kQcRdf4dbNl0dt7uF8C8hT37nncq2
mtUuMYTtQmPGq6JE3/lV2kKySlZA2dDr0xM4b4L2d01OVGOm7FIWiQLDt2oC0SYX
E4EhYQaaAqrj5tFknEdoFDuxFelPCMaxX72FuIefVXooOGuSCMollg1cj3vHI6GF
L0FBgAyJhM+wqjA4ldiRoR0922a7qjGMFn/yFZbhQepLwGKrt1j3wVQCL2dauk+p
RiakN1DLIx5u+ZvapXtQ2KWh3diwCOYiQBT4uqKLfscsEiRoM1o29A8GGpc+X3Ib
4Cenb8I6IkIXsJil1A1Um+lLpHH4P3JKAzbCQjq+Ks0Zgew4JwyvC3Uxno6M4HeN
hiD14IIY3WMCReE4YcSHJSZ6X+RDBF2ExW5/P6b9rk3MnWQNgq73p2MmEW3EZE3z
NK7gXM3ZYeB3oPhfccdhXWwoeSm/Sa0vVR5XE5XXNtXvvxIuyz3JTPvMSOz6YWXI
OXXvIyZD/5RtEpYSLJhQwbp1Cvgq+WaNImmJyCgXEeOZIcVfi+SuVye0kiYiW9dm
nERDG/yeaAi8yzko/lwDRXId3m4loz+4Z9ZAWxXFHu76rp94nPvgwpLBzHLgKjKV
k0gv7xrHYQzNs5A6lEp5f4YyoerhJZunsb/+ARyq6We++GTsKBMr75XKXFR4t+Ie
fgnJaXfsHxnlmSx8dGqb6ulpufdsNbIZL0aPoWjaGubRBamnl6objyAHpmuk1Cqc
ndrk+9RFhq25e8FPlpBZBDpqdzR/s0SpoS+whlXx7DH9OMKJEM9C8yP3lYRGrhAh
dpigbJMugh9viiz8okyyuHLTAtBuP3gy8piV3vbcaVjrNb8PZS9HLguRbJj0ZISw
FyUU1Gv28/xh4GUOoNi/1pStzwxDfu6zFWS9ocsB4uLYGUop0dOziA3e/SMnSgQa
5AokTnkjKkn+ScuNcxmfC2bFcYmL3cwovSkjXTe9lay7aVjiUUZ6pqPKSaL56jIL
+nHjnAFAd6mmHkQ8DMKdPKbOapVDPmjiHLNQcLv0Gvv9Pp5fiJrv04Txu3Motq+w
QbiKEgYwi+xdzUbq+5ySFbpdXXKyk2xrxomaCz70AEB+EkDrPAVb2UygFoiEfTgG
Q7nF/OOpuZfUuUqBrb8LQYunE9p/jdkyF52kQeADHuMdE/aRGxwRpWgC4Z/QLTve
+UfqCTTFPa9JygTq6/0vP41u0INfr4ttMStUlJZ6xg0pNY3XrGffHb1GyEm4rGoz
ZK8O2PubfxJjnK/sqJr0Y1ZMEIBoGN5L/m+AhgnfflkpAyIxFvnlYVHCIBhXJl0W
npr5WKdNc8XuIw1GvXqVWNY3K3KWf7LeCzY8+bG7RJMgH6Pxb+jX15qMms7vJBdK
RCAl8GKBV0e26HLxAEI4dt21Z+ztZNumLjqpsETFJWJIXklMQ9tujUmfUAKCYMuh
FbSgz9DUtA64MM6PJmIBPO1TsvNrra2XV3VSVkh5EgsS05kOgrvxXV2SlQn4CPhV
EUpeRw2DUnpmU7IN90Q3bqp60AxuvxvWTC255W013AzO07dtydJGDZ5A9C3RLM9q
k5zsWMz4reAIZkiXu7lkat4lKHk0p1UtudoifwYt7zsteGK070AxWyeCM8jDfL12
0EDcP8nY7gj29g9cU7f9Z8XyOD7rLf8F8wvFfbVOAvDQT6RaohdvfHbAVkaoJTG2
rCBWukeLqPkgw2p2oUk9zEgvaLYGvajgJFAPIDQvAkqXWulby9SBTAoHSLA6KhWS
dtNokyJ5/o88E52ETfo6eNK19l0GKqgkMl6WCvy61tWWe+SVNJtwi/YB2T/jfq8+
G5JfyjAtYJCJ1zQD73zIGPefY8+05K4/5etBRFdipZAsLsg+ph0K4jG/aroqQHQ+
N8rTJZF5IRRPK8NvzH9nYQWKWPAM6qqFdEVtOdkE0fdoBmjC8JTZ42II/7oGbA3M
lMkB52b+uateC0ovdr4J/7GPRMptVO6vh21bLaNaUiC4+X694+0OsWJpGzWpFm7l
O9usOq1BXKp05TIcFH8/FIGTpHhnyFEJYu0wlKrJqlcfUkHMyoINExta3Pp6iGjP
7aVTAvprk/dqL4Za3RDe8ld8L+J5Rj70QVC5DNdmWk1NEfaUh817ZJcrE5rkE2Jq
9SluHJxOFrAWS8HtpeE//BK2syE3JE7sjtniUukZL9atfJ/AbQHIpH8MRfCoEwTl
McCTpEujhu+216uE2ywLW3MAsxpZAN9n/igevB152D3pJsiREihlxjOamJaCu0t2
WSu4fNdfWtMMhCTjYGxO5uOIiY8WNR+/412bg5tzqGdh/+C06PliJRJ3FE/5sq+A
eNKZbFv1HZGCoLO4aRqMkj1YwSgzkjECO3vBIv9NCm1JQZU1oWLYADiOWIKgh+Kn
WMv6uAVtxF9k+azDOSPD8lpMwcP+NC6w00QiNbOLY7PrbLYpeOKOvMOVw/ezwed3
t+RWFmedtiR3hXAO9ZOjD3ca6DH9q+8KlpADa8O7TJwry+bqB+T8kKi0EoPDUKiW
opn0eYqsnDSwfPoWonLVyMW3fXsWcOQhqys82cAkNX/+3FvWjID9MSqPUOjMmsZd
0EFl0tcPlcDI1uBQWtanYJc12954bjb4Mmxa+UDKiA80+1Mf7RDsf8boqy3ztPzS
E+FR6EdNOKHNSkGD/QkjoCRbRODUVnD/fxDiNZoBdy+JJxFLasW8V5gVLGYS8m1M
+myH5bttGWHNc6b0J/CA/Hq8m9zS8QZ1Ul7vtQKbu9Y95nHzhFcYVavPNzhomoiU
NO6r71CIEeEOFTeWXWmHIfX2mKVhBeOHfa+L06ZCkh3iOiBvXMBwhnPcdkbFNtrf
dkZH/GFZ3FZFC5oFn+Sc4nomd7hH3BGdjmOFLt1FuVuq3dl4EkFGuf/OwsEtIPbm
08N9nD3Ia+ScfgoGe6I6WWvzlNwCbPW7VkYuVfHs+aJ6Jewj/UxPUIyFK04N/eyB
b+JrJ0XUsPg+RW+FoyKINv9DBFbsPmn8XfBmruY9+TwuNKB+Q+a4oBArMLDdvraT
idgtFCgqSiZHEW3LSVRp2LXETs6Sgs+jTWItICG4v4vB8R8AxD874Wna+uE59e7E
0ZLF9GUmFD1U8sgnO9/uqhu5nuZ9a25OlKg+YlfNjxMYO1XQ8qY701DK0vb465gB
tcU8jFzPZDX8RwR+vKaKos+WSD7zriY6PDXxUuaWSqVgYnFbOsuQA0qeH3H2lADn
o5UsvIJoJThMn1EUiAFJU/PzZBwhT3UNFNYt74KEQGZoKLA+qSNl+8haRqT6XmcS
XVcUpU4Qft90wlx/WcrPnIWfHscBUK7NVw8F0wQ+C5B4a0zOuXxVIYohLa6MhdYg
YATsx7Z3gbCRKBM4OLhY15CXAYta0VUPQtyU9Tx98ooIiytTR/l50MSPLG7fNxye
ucMiZ2kCqsa7jxXpQc7EHV80ScwS0yOp/Lq7MV1Nf3WMeB7ZxCe5pNCpdh/L1Gyn
tYRy4c9Zf/s7gmGvQLURbixgqcISyRIyciNHiSX5Tb52jC2H+k2F9nG5rrWaTE6O
bFjo2oi9wcSrqRlX+dkEJOndM0Sop+Z5Dt3lfqFUYJuFSBs7r3nkb+wHjMtG7lue
u6ALmB58o1s50Ewtu3RT86tEbrxOIJEbe6Oamom0a0omueqgeKldNVnJxZnJ2pRZ
Mhaj55P1GQFqt6svZ8Lxc7MjUVd0X78XPNUU1+diwTjF81YEiqQouajck90wIpPw
WoUtdD5Amr0Nre3KziYRAN6sRgjqn1u3oAbkWimIm49GolgXwMbO5ZwelvDYDV2W
83ZDF+nrawUiZLf2GlYpzIhkBSyAXWXVJQdnsjQfNc43e/uBiIHoYp2r+kBb3kWM
jePrO8VOGUXPrQixwCPIFmt39erUNeWXP+2dh8zLBzt410W8MgQV8f+PWr1xlLkL
GmiWfqp0Vc6KAF/FT7lizzro5zEVk07PzPJmUXvB5KZLAst0atNV70KGbsqCm0Ku
5iBdEQBtJY7sAX/Rv642P8SEs4STEGDL73wTboEjwLj9LWxM7TNlcCK4MTVfP6Av
gxWCDNiSZM/o8JcFu830qnpekO7zo09P6QfI1pcFdJvixvzL9rXjQaIdAZLFR3qM
3dlNzvHMMWS77vveKuCM0y8PGqbJpL52M6gzxDKjXVhLIDmV22bnMu+btlHf5dTH
zxki3CJcKBfBBPdUF5limBqZQqqCobaWHrjF0fhlTIlu3Tc1y4JraoKMRTRQm5v2
7heEfwRfoc3cdFInRTxUjATC7Gf6adVzmOCk0nOw37GCspZKrCmO/JYD0TMQyrZ0
sHPJDsZXnfJdfb0XBkA7PE9TZZBe05Lr0hGwMtNknTqamxWfVk7L1YGAt8N9gIEI
u87i9NbnjyMaPml99vz0x2ofvHY43na+h+WY8DUjs8tnZCt6KXOe6euAgoq6cV+x
JyVzWK0mnpc6I+35HE4CLe1ht/HhVN5hQAQuFyXrW8kg+4w0+fNdSS/7JcWdOVxV
JE1zbRUJW7UjJ7sd8/570trahSpzzPnCG19nwQx4lOkC8dOfTYl7SjJGiDyo2luo
u4/YtqRlDrz80OW7Wahc0TA/H+qXSIwpeajF57/J8KMls40npSpE3/NrjdNLwO5B
0TABL1GwX+ck0BAX4GStb/djBALUglYjiDTkQPw225cbVzV3u9MvGHT6UnrdZcbf
+b8AUFeynmqaAOLaSDCDu0lC0Z+Rl0FejWAno4iQ//fc8pBzEEqE+unR8EJeCAYH
JEJGr1AfUqDNX78MAZcbmZhfkN37GyDVRc5cL2d6IzJQoFINWZ7Oz7BWrwk/XMR5
vG0BrBTr+52V2DY9zx6ItvOluGxZkHvF2yGqplF+hwclP8t1VJ9zcT6hJ95OOUZf
Sb79/E0SS5z321PAA1sMCWo/iWMFrkD3UE12vfC0AARS9MVcVKnQk3cjxOzOiN9B
8L154iMi3Cv4Bdd+anOr4KoVEbiZu3O5fqjb8sc/EngasMQGt1e1rxpOi6OyDvPC
F90cMcmZdHs3JT0ikJIHKPv8lQQoFegpHjQOo8ghg66zNaF78VICa177I3mtdUGZ
eXr1shMYPVnravNhSX6YkVdUuEZpAvwAK7pcfh64SB9elp5GCURoOuZCnB+WSou8
RD+GBQYDw9yQ5MK5uqIhOIrddPmlb0hPrzOdqJgfoBevd2PZPLDKMSsrJwEA6lI8
f85VaWfKJs9ky/HdTEOPH1CVmOjOVOYrTkMJbCGTqBsG2/N/0IF9lhTBOVgpAVfQ
oprXbLhODaDe8WHnvSDcH20+1NKU8A+sMHRn0ypTCdEhyQYOJD0GT+pTorYlNIc+
qe5iAjNnaoL2/8m15CDtc9XP9W3VNZ0zhoBrSqZWTFHkqsQ9/JeyJ8heuqII8JIA
wrgBa32xkkThLGJBRcrxIk4b9YNGS9myeS4UrOE95uBC03xGghQfZyEdlv3KrArq
e96D7tXsaF8mN6PJSSsKr8iH0XC9GCkZn3KoIbO0Wz/2M3zrqBwE/k/yBnzigWDy
hBsyG0ONe6ljwVA6zxpkwvr82lmHsS4MqI7lZS/+I0XwIgnewraPGNevPy8GdD75
3RKskAha79dtb/bEm28KnJ+DfdfarO9ShRXQfR3x/vdOsYM+3VZea14KKtyCOAYv
9u3cbBURaJkwxtiXLZwzAfQAuzYc7pWhpIOZNlRFTui6Y9BHoogUtUqlkHvHXvuj
IsJiEzhxyEQ6qYZTsm35Ge4QebFqOTxik49iewyMRdsDzZxJACJeJSYyockVNXOJ
VeDsvy2KAW6yc13CAIzrWx3jOWtraIWCL8vI+xYXC6dffcnqURXxfIawQmOHndKa
AEed9XPoS45Dhdhz9zUbP8cOyC1qKYbwPvCWB6OOxu/Uy2ffnszHxjr+NJkgFVim
ijUch0/EcMnAVgx32mvxrnHd/glHfd0fi5EYpQ+BNDAMZceUbYbAkGZezIuP7Xu9
//xzqnyGVFuBcWrr8jdo7aPxMqGyrAybM8UkiRNysOQC0KN4Pg9yvOs8flqaG0f4
tGtAwPzt4ojlHMsQvHjnYv2La/ld6hRAUX/KsYbQDGo3JFE48Ky9ebne9HENO/3l
Odm+730hTX/NQ+3xR+6Z7UwxGY8au7j/dQV0/eHPlw7x97fmE5NsLMdhttz1WsV5
NHMaQqCwmyMdxfkWJ7uRshj0K4/a54NUR+hAEsWqP9keROAGoB7frq22FPfPqPhg
pOWhBD2nSZfqOoVVvEXVOhSSp2EsjneIF30iBcFGLe5XaPq6wZi6lOG26VPnFyNw
fvTD4VmQGDpQPaKT7KbA61Wlp5Uaig8PqCgIgb0K7j+tDuF2pingABeqBozgV+gb
WcQ9pJmcHL9ax3ae2ix3o/i3BCkHi6tJK+8vSs/cgq7NqQi6exV4jIUWdIDlLgfY
kAkUNoR8bQXiRN0x52lEI/T39YI7Q2P/9MxY1hPt6yRY1kbIdUuUswiRQkiYitiR
VUrUif0WzLQuV1hb98S7D60OmVXnaBSug9e7SLfQFEy23Gts6ZOIvEeu2K42jPqr
sxXjiEOAPkjNMsNgIYUPMjLvmWwj2j3Rkjqa9HUqLRHMXAK8cKJfE4JlRIn+kqBc
/O7/tkLcjrGQtIVp5T783vMOGVcWXFd6/ko+le8Ot0JN6UCxXKDThR2Vz6wfc562
ipxhur08SZU5DIqMBfwkC+k0SI3twItE+cAv+Su/882aXtOFzCcCveIkh/RARogr
OxHnUMYL6ehDkyqRV2QZzXsuGLr7prVB7PfZOvFlLLh0MaK/sW0ZPPBRdLZYMzcC
jyrprdu0MhUc77hiX6RgyUQLhmvetriUc78/vF8POn6McpeDkPat99wdYomO1mYR
w9gPw4lPtKZAjEOCt/SwtlsLlgMWtQMtPRmWWXqxbs73mh7rH89dxgf+R8XHhTVA
RzoZMZd69JkMcZRpCOrm94FSp4YCKN/8P7me0eXUmakwSZB+tyojl0xRBwhZ9diJ
0K6StBrXX5W6wbMoEDlxmobsy8+oKkGbLwE6augO8IV3KuDcrvYnMTQHDu5cUeOs
5zxyWnIeRspMaPvE4xvMKkxbzf8AT4u2qEKBdgyedhzt4Y5eyeXtbbKah5TJG4vO
HVzh3zn/8O7T281oZzqaTbkhxbOy/Xd9WXbG+y8TGwSRKezZMq8EtsFTPBumK9CY
7jMmNJuxVwgLaKCpiXGz5ot7TK0jvoqGBzVBHAEeZd8Arzyta0mLft4/eZbMqQL2
I5CzpWILZZk9ktwnEIPH2RKcDUKlPKIe67pia8BCpOlgbP2VZ5TpsiKZh7afgR+l
QFmgBiNxAm0zAiAWd18xbm7tqS3CxI5UURDOoyUmlS/7L94r758tw/c8zR/z3Oq2
iS7l7aza9FB5bSEcKCZvIkxuHm0GNqLiJIIdwLWaujYZtj5r75DtacB7l2IbGyH4
N9iEcB/SR6Por5wWOow3p953RWTPuxJkrNqPUOXPktM5AO9tKTySsYQUC+PzqtTd
5rYvbM2/yOL4vayzZPJ2d1/XRdAmlXAYABCXDIbEf3cGQHO8YuAVQplrKIl5wt/D
6Gxw+Q4D2FKy1iZK1l+KylQHy2XmVL2kzLTdq5GEjNdJBv1N+gEvNLTpvGdyCbSm
N9ChfPiFDIvKxhWghKtWywWnlezA93iLzfTLocc+dvnD4y4TWldcQVUW1ngk05GT
MdC65dVJXY+z6wgfQYRLZeTnZUKKc3E3GN2fFhJpnAfmNoecEYd5j0jBlbgbi9Gd
bKwtyFMoJXVHieZ47XCfNVeyKXQWDEiIokr0xsrJl88VGZT1ibk96jPU8BSJoCUs
5ga+GOE2wif/8yTiKdfJNYUcQ82BO1CtvSFMe1nF4YiaSaLFppmWOcEgQhrXmTTY
6QoE++i79FpuOAFoAGwhpD3LU1OoxfJeCwziZqRt8EEF7N83uEnsUodKqAsM19sy
7gjeUBojxX+xf5rewknFmKK0olCPyg8drPu24woL289r2PaIN/GfT89zwH4cuMY/
nPXUPRQnoDALu730VrntNaKsHMGW6M5LEArw3M5bN4SzCS0U48jhmWzRv+nYGXIy
kL8BJWOjfxwAdTt+HFDxdKpYs7w1S9PgE653+3C8sPHP5yg0/1Z0iKf2D7ACtFAf
/ZZkv7xh35OmT6N//Ryrq8Dr6b24uHZvbGkqiWk77GrY6zSASBzQNOQALEqQhtIS
9BaCF72dXl3xiRR+R4I5JFa5uXMt5X6oe1KFECq0UrnPj4HyUHx9RNllghaV7uKE
1cKmwhRb7/RFVX1GoNE74h93OS5Ggwgpo3yCkt/3b6cEMTuR/OpZH/JkAp3RLtMF
FVWepvr4rdoHqr0q+zZhM31nntBLW8RLP60W5Cxb2eK9pnZZF2tAFjO/uGG8R66U
9XNfA8UyaNq8Qi3sj6Kc/ok/bYqVpVZvx+TlUT75J6Ji86e5JdExv2JOhtJsPDHq
416+HZb4xsF49KEjvFdnzojJD8GseAaTkuuCRLAqflNm01eaF60z5ah0KmLWuNZL
MMLlK9Q9tZXifLM0x7hL/JPJt8aiLRtdENhcDhwwcQTKzUr0Y/lHotxVo1NQ8S9Q
EQLNRPmks9I6rd+i8mc53M7YLGN8+Th8W3yxJPEgCibLyjslbCMBAINDVUr+37bF
7tRIpQN7+Q+faRjQoLcNZ+DtGBqHqaHhYFSiU+AadFRHSVcHUncLw310wQnBCheP
4k08sCeOqaFsw+641qBzK1edLFwPXWa5HD9IXHDR4w1yGr+XXnT+TRgkaoqFk0de
mEwDJwlA/7pHb6s/X81CiOL+8WPtwhmoevqYVwbqt29olijZWWWwYQl3Ox98EkA8
U3Jz7Nhy9zo9hUUDkS3gOMYLVJ0r1i/KM/twqw9vVdLgkDtOSwdS2LcHDvdrvyip
xC/wg8PrtpT+wqfmEMBUNhGAlYExcrnVrDPyKRVPH2lGFu6sY95KRKjEU9+Vrhqf
hC1U0c4VTwCpIphhIyVwLUcVDTsjDycjJ5W92UDSx+N3drnTBUxR9OA44Ui/5c9i
3sJwvRP3rhEDLBn4Hqosn2GlcqLEGElhg3aX71fVfGus3jUrQ+N3AhVAe9LjBCcL
ASIMCqe6R09NhNd/BtqyHC+b8fIml/bcePoAPokHDVUbky0zj6QTaTGOICJqCJyl
eeSY9/Tums+xksALnzk/+NhkRweGJX/+wzBUtfB/a30sPxFeMMfOmU1Gu96TZ2eW
npHwtHyqdEgGsA6p0x6+XIFLZXpUe8NKn9gc/fRJlWihRRw2doP/ZwKQWNrGsi3K
TKJ6f6CerFiKTExh4r/LDifwGxcmGpmqO/rHYBn0YSYL/h94I1hvLZ0VNVlZX45v
o6k8gwnOJsJeQuX1pkz9IGXq/s/4gqReQHyyVYS5lq95/INsk7G0ONfslrh+15DZ
+rBX2ticSMtSXVCNivkhGPeW4VjARELOMHlkLdtcqglgI6yRf0GJwe8hkUvG9WAK
cj6mZpgCx0Fj5b08wxEZTZ6oF+ZxF/9YbdL4F4oOhDVOksemp1ARBJ5oV4wUlgQc
kdzcJZ556BWu0cxDi50p4WKMh9omGoK5b6Iwp2WYHb+GXmi76FIKtYjRDCR6KPgA
JLDdBmkWzfxxEOLtwu7Fq0gJivB7kqNzJdMOzbd4xVnOF2abKDUJak1Fcz3HA5tJ
xQxfLenJMKO26FxpLaPabC7cz/SsVeqIKeutbEaG7uaw+cS3DVfrYIgeRnW27NZ9
/4hqepL0ZGyDxrvX4wZF35ZfQ4YLTidfLRWFgBsjyCop/wgfl8ct74xbo4d4lc1P
44G2zXjHNBsVIDbo8U2UD7UnO9ksE/T0k65QjZXyLKTAwc2YlLtdZlcNxoWTkP2K
PrfHYqQvNBn5OCz5XgTtN/FEkXPxVSSc1MFVcBmX0Xd+/RepJBRT2kCZkgI/OO7r
U3L8n9Vewt9IEaFc3wnqZtMhbfafVBGYTU5eIs821so1X+bQ/bBaSXT/yezLQj83
5MUxAbDiatJMxGBKVZoBq83kQmHsN6aks97HSLfepCcmFNO1Bpb4NluRB/kv+ktC
JPR5aHTK1L2O412p2fwiE9NOInDI7mrFcLBrcmiSXB/bIE40EhT/2SCDg+/mek3u
QkTbkf4HmtFstWsVYXUKZ6+PF5QnXEc9fZAIMFdk3iKTcRh1xrHiVMDaURpu3BVj
+C/EKwzwY09W9TSWBP7XFJN3/A0PzjnzkkNx1hk/UGf35F152nBrtCUBu+QF/hcM
Hs7Zsv5k8XWV2hYLdRzCFJlpaSIAVkSsbojM2ZwlgwHyDnNkSXjub4NL6BPMA7BI
pVCYuCJ7RPyXqUZs93N51o3M5asvLKbY/w46h9ganClKT9EPE8eZ3eMAkmqjHJ4B
VPplw1RVW6OxIMBMve2P4HRYI8Iy2eQWcwOdp5nE/j+VvhDmN00z0Hsr5CLUgzNB
rkmRgtwNDLyRbVleQtelZp0D8Z1tHdpSTMIndydYi6UQG/WChJ62z0ZJARK/Bk6h
Zrkftbn650Z0qmclBrToonKg2W4Yh2qtQb1GXxlWJF7TnRIVEcBrlRFeTHuTT5bZ
VvW4JEVq3wk4JFkcBnHmwUru5hYoCcq6nX3H0j87/TYT6ixqgivv9kHo2908DKZP
xx28EpIwzRIlZ6hVms4R4F4DXVdZW5eTj1VI9JLy+iycaKcwf0AuQvRdWWn12kFP
BmP9LwHIW5FKxYWmuneDzarkglgrHA/J2ezCamixA//CuUMGL/NAv6uBN6wKTVBO
+6Otl2+KM7jLKT2+sR4XY00Oj1Y9bWEcN9Yd1wZb17/Xa0u2/2KjwqZR0B7edGQ9
0WZQuNzMZ/FwYXEUw1U9m5E0cAzVubhnOH8cmLblHN01Fm02vwiCRUh508Yo9sYn
R8QPZOE11NjlmNLbx76PrD6b4Ks2y0zM0ijKKazmN/GaiikLmmfub3J0Brd8l3be
D8IscMpUxCVvS0CgWZnkqIoG48hSs1pQ4Pudeg5lnEtURHRqqogBB7cKdP18eqet
Fioul+YZM2MKyOBqCoXiAdDqWDBnMrvO7ZZhHrlH4wZmlqm33j4LklLuFEkqxKJG
tCXVvzOlNjLmrk36RUeoDvmhJyMLXmLpufRVm/mXp6IVlLuZEijzoF1NV1EB/6SO
j02PAx3TwvDOQPDuRwSMkDlZPOJRbkAu9p2bbyt5UrCIBwyhJsY9r5JMl0hBmsiv
r5LUVQQgxNZVfjLmFgs9qYQwzLfZSN9hqMJNC5mZVqIYpBAegbyI22RTYePqJxcI
1Rsq3c7oEalz3cfy6rooGHSs292dxI2dDahLcPS79DFcJ/LQoXVANI0FTJ2z12/q
PlYnAHi/2yA41RGTE3ai2bnzzmnbG4ki9jtlfy08xpqlqY7fvepQ3Ujoj+WEmvxS
KO2ExJkBaoPPVq0zbZqqO39em3GeoN0mZdiWk/NITkCdCAfTTT4ZUAy7WVwE4bOZ
nfoectCaaCXdaLk3zOMNqjm6j/y9ZEyA1zDGIIoLC2JKPiNG86uUOYoOhg7kB4fi
OUWtX0ud7/Qzntr4K/YDEZtwjCMpj2HyqwYubcIWP28CkXdHgSPmAmyzypU7R2ZN
NxIpCdpw6jEfkdelmvNGMDs2w/tIAnfCgdomlm/26pKkzNr/RYPLa0C74Eifywcl
lnR1Zn/pmhJc2KzLhf2rcrV1QQideSNrztl1EInBvC34hC8N68DmU+QXjUvZcR5x
qRh/MW3IDiidCjfQvenSFIZpHL8fFineuJFwQgj8EoX2BOwCGwzm4Zx8ab4WK3nE
HheKlD+SXlnQY9G0CuYfExzz01G1iONfXGdW8DTRnRNev77YkTAWlXJOoQ/BtQmE
tWquxLQ1IUm811R+39gGcwc9HnepWkKl7A3lJDAyk/nleioo83P9gdE3WV3yFggE
QrN1NOU3AcIRH/PrAy23LTBLRQ1dAjJU/2teaF94ouslvC89flUR8TRA8UoTUmL+
ZdKAtwCgZaUXfk6HN3TboQZ26p3YWx1Nhr0JvLSYBSD7SluNrjPN2/cYbxCDxsYK
I+BbGtHu+4QdSycvMVWsCLWtjwn7zbXeUCsDSFo3TMNmCjGlhgDxePV+iyTPY6xn
vk7OmS6UdlT8TP/NZzQjGezuJburUzMngl1bg2WlUwhWRm4nFnxPko9ZRIZaAOcb
XGgXIm1ge6uuXR0F3a/N03cfEcMbmSAChPouaKEEwwc9OySSn/LDeQmxWdnRlVEG
6pIi2KHVnQfBsVBqpZJrU5IwtL0VLQ7Fgq/JcueoJnl6pIM39pgx3XZizJeZMkfK
i4AYyx9bjSZfIqoc6w0syK30vmZg0/rBL7N304wn0WVc8SJqMMTJf+mEgQdmYe3e
ro5qYy0n16UC5Hn40ZFw2liwnAC3DX0kD3KePSXVjv8QziK+fpu6Mwc5k4oETbl5
ceEQKlekxsvYyIJ0aIN06nTNPhovE3MV5ifdc1og2oV1SHD/uhyM7pY5i1njQxoX
oo9KHkcA2ttxu0lkI8Gr98ARc1jRN4E1v9gzjmxaizUBFUTWtOvQH083zquwGshd
STqkBWXppz3JtZo5TYtLWaFTicUg2y6gnNw7wuzMIp/z7pX8mZKn2Vy9jxWylKf9
yzJA69XLJBRxhIcUEeYxW/X1JrKUd/aIIjt1CB92XFdVQk0p4nNPpQrbslETMUHb
ZcFH4eIaxZ6x6Y0H3rCwzI/0BHwkOaoKe+uHpZeQogwmBP0SmYGKfpbtA91FRB8C
LfLd9a5eMnWPsbyU/UNGYpoIbCZHPJvqeI9RPhmCFHLEU/7Wf8W3pUMqe+W9dJRS
CcpbQurN844lZP5rB3JvpM47YztGGaG5EZjvg0432/eWKHQhMz8w9Az85YZWQ0fv
hCg/Kv4ew0xT9aVnFGXK8P/iYpKbOjHqs738vuZU+3ok5rekPT2PHdpzaxMeH3Ma
UaW7pbq+6hYBP6G8GCOMyMCuUCd5P822oLlEcDoMCMEra5s80U/sTRSACJzlWhJ+
3Fszx0eD7hSl8eOtf3N6VqHW2CYL4t6TgNHkB4suvsxhweR/vhtCp+WC1wPV0nB0
M4kU1gy2VaZxlkVVRb3putupcOsDIDVpKzqa+2xQ1eT4/HgRt6DveqpmYykr4sXA
pDGvWORALotsuEh39o6vN1YgZui6ikP5n6o4QY4qpYFLpD1J4xw+p61HMnppfT1r
3u49lf/dTpusGL2YbMo+gc7DGV+W2niXR+U0b58IsWmEdYSrTjiykcZuGnMQE+eo
2NXP5oMEUrre2yPhe2vB1h9qXJAFEof5DNL/L4JlKvAtMjRbzMtxqCWx8CuvQ7F7
gAptpvmzF0lT9O+Pq+AMVIOA/FpJpTg9IPQdoqLJFH4VQFyFmN4sPSh7Ld27sK5p
mWPUkud0jUXTZifxqt5+eU01L53IzOuDB8rqTNDy6A8iCeAMPsNYmFSJnr0fcK7h
UsR4e3QZTyorncyX9TB/CUEi2VYzDvWLxT6p+HMzmdm3LjQ7doAHBfohOoN+4fDu
Y3JGYAmv93ks+iz2B4AkLppdi1IKtqbx64h9RymAnOARAFu9TT53ULhjEuwHTTmc
/L5FwNq1/MYAGhA94fAfXcTzv0MUl6LkDtgvbaL1+PSNYA8vDy5gWmwduMmnWVAE
Mni4O4Q57POtS3ta9yV8PujUSD9q6ngdWCBbv9ClHDh0gr9QyMDEnk82j/Jyp91+
yqFJADwFnonxMYLSGj6blcM9OOgvWxLfCmkCv1W9hsdcI2wTJN3LP6IDEi6Cr2bd
XtVpKL/Dk+6enhifuJ0eakx6Mdt2BUJVyVXoR9K2EQ1Othih6u6l+kcbvngZBsyg
jztDXP9JNYcSQqXb9bjhs6k3AljNyTk88tMG5X/X8pl4hZjkXjEvikpvRg06aReY
XGJAzRM/qKI3Br3exvc2S9GGF5rBzeIGL53gR5LfFn4qUYQ+nFcaPVnmzpw6IBfs
tesAYBJSwWj4xBlL5c8hcn0j/Zc4l/UJskgE2C9ZsJc9vIaRRtm1hpxMFkmsuNXV
RwZQteCC0OvghI4OlTCx+7Yo8+455PBcBQXvDs7noo7BnZYhewuxtvnjUrLyqYC7
BalbKCvJnO2HmLaf42MK0ppG8xTKnzdqv3arOAV+Z7Kvz0QRN/wkqZy1vdjSzwE0
8R17lg4HmaKrQvBpjuPZ5mgpJ9X8LEVMG/hWIXPpU9BlrNRggSPcHuarLYsvoNxs
cqBCtjyHwkTyO06o1fMIHikHykuu+C2qkJqbI6wtK9/uqekU8T0BQMQc5Re0MLIS
CFOHxiY7xrSAlmz5RlTNA6/lvaea8J3WD/RgmC5cT2BF2FfShiPikJkZCE3oHYIs
MefjHu3kDL4FHJ45U3DfyP2ipKrEYjOlKLLzqj7IiKrSkA/v6no/lrcoJiucrzT5
d4oiUkUaBsTyjDnEDGkWht7U+/RU6J+SAgWzWVMWh6wa2j2JfxhmPqMicMXvLa6a
WaB4iWV11sW7+CdKUHenttQeUwv5ZKvzu94RCQRk030wcW37M4RBGBPQmkkyKCSu
Lb2DQAry57fAcCkHWZlA28o7yc+des43Xabkst6WrItsbABh4C/eWedmpFq6VWfV
DiGYllXCSDQD1qflvKq3UHMg/vVEOk2Xb6rZEDuOooV26iDRoyd/3TBTQm5tl2tb
S25f0uSevQQP9ypk67FQZqs2aYxrmZyH1ueAs72/Ks8oHDIKAFXFQB8npf/L9IMK
LxzQULd1dbXvYw5BSn/DwfMl1kfI/BIwDA/XWWsAGPirMoohrp0O1KiEct6swssG
bNCVdnrZ1423Ok7WVQ0QviJPpnkFHmvUJcC7pq1nnTMnw165SYUIzeTPhX1gkRYs
aFOIm1tadvBq3N4sFY2Gc93minECoS26anrT4M4m2dIDQ4Z6ghpOzcRn1pM3kXtH
idxxFnEvBOPULs3L8EbrbKFFU3fBjggm8STYuvCyilo8+ZD8KIi+fi3fDtzlkVdh
gMdoV5fiamhyvenl/Apmrmlx6OhAuBBcpAbYWQLGbK0d5xL6s6GxwtSetxhCWe1b
ZhVSbxxrAnm1NrB2Ow2K/EWeMbUZH6s1efcYSQ2euYCvOuMYjETCnkq7MVWBJCYv
R0xeOVWE8rzAHr6exdeK5yPjumLY1XDb8Lppf4y6dDyfK/z0KURktYbcqOK5m9OY
A+7pvA7SRv8gYvDEc/eXjDNGSWmJZKVJriT3OF/2jwEOzG3eT6NLx4FymVandvW4
EAwPdbbC0XplbDPHyw0wC0amZiDFGoMs/PsaapigUtk/cWMwwY8U3R7UCyzi4uFx
WrAT67xv1tIm/8B9QHAN63KqySE+Uetk19qkUK1ihczU6soav52Nb8VlW3rXAo6+
HStbNHvjyQ5Cy0ZIZ94/9ejEsFMI5d5esyOjYh0vdMzc4zgxVxRJhelbroHq91f4
iwxplLFmLXjpQeYiHlibj1Nr0ihskoJm5cdRu+/jgypKvXoPb7bBN9O6WmY6Lf2m
0jJ7p5+1Ps2bw0Jnto6a3CMguEjIBM9pljaZkBk5UZSXrVZdLPquos6Jj3H/w0S4
LIgAvGuibSNfq0tkGTNKB7VwY5vTTWANnVIU/vELoOjgmZ2dH7CaGHw8wAzhWk0N
aqTAXmJGEWtyr56btNprx2uu3XpcOkxuqN6WfMHbq1W1gQL0RYNrzRoRJACbpvUd
QoUbQ84MZjrt3anGns8hsXO6vK/CEsxxGdDYqMj2jrI4rblbvtTkF1y6rcWKQGmN
H6XI3om/BqOG03qhV+4HtBTlnWDxqvuum4VhcxTCMTjrayKsfXnRas/8+XUV6Yh0
hA2VlEFmBYPIWif2OEjx5sWsezksXwt3xLlm4Jp9tXbRDe5b8txprUemWeIiMSMb
xBNd7TSk3t3GpFqWJ18IOXn1CZM2HFJnhD3YoClzN9bTFmuTveWmCOhVg61b3Dvt
D/+kqAnWjcBwBRRKGtAn8nn0B0dq5eIvhfDzf/yJXd8fC0ojlWRSIDWnE7Bdz67J
UhGzMPkmnEVhAtyUcUgZEtf1InQrUj2ZGV/UuZVdiNXaQR1oZ+mnFZ9fEfPh1TCv
0qAxLDbviJ2q27WYsYQRVOK1/QwzyIBBYIWouWqD4D/ybYZQN7jiiO21Kfq5xxC9
0ZHZAnTkhaqnGZejBxCl+BxAdYUp+JIq+/Wi/9aY99v9juOf4p1mXUNWrEf2+T6P
O/JHvIU7a+QuNmqPc6ad7DOicXg53Wh+aJ+708yT8gMIzGvjkT3/rWh85VSDUGbv
zTxKhOMZnSfnchJti7pwYFn5wy3svzhlBGqC1OlMNSixhNVYQxKxLS/asIDjuxTp
IgcAF54Fq7LC7q394/GaIs4frFgUKsL2qNzl5JJwhPZW/W3CxPf0VxVC/sXIUxS0
wYUlnurUeCApOdA/Zr3wTbdR2jYEoV/ob5rEjyRQTr6at+QtjsEsB2+iIxnXX3Qd
hiP+qs9x52TziI45BF/GUdBdm/J0oTwzqE7aJ0EiET7g4N0J3zFAk7BSVp0ke8Dz
b4/n4DZtj0YozvRONjcj/JvL+eyxLeBaBCU4uhPCJi+Dy+etlMFVhEZQJI1EZvTo
xRReZ1obI09+MNwN9uP07mxhjDS73p79WerjPgyhY5Tr1jz2Jais+iaWblupJ5od
6jXX+OVu/8riyAnQO1pFMk2zv4H1f4tdBpO9rVoCVhFecgXsLfbu255EPLr2b8F0
Y0xKWh1GBKKKi3s8ydNo4IaEYSxVyDs3gQx5y50cRxeoHRXn5/EONFtEhF/UpSxU
c4/kZ/hwFxIHBFAB75QKtyVdHnJCP0W+mmZsHX1DfUwk9qfHnFx3ruiorQ23FG5A
yOsjc5KNrrtUP1q4TJli/cr1S0yoy5g7FgRoE149X2YbwCCCVpO+NBBLDomKi/zu
HhrNkmUxdnsU1ODhFD2dvBJXprL+d6bFq5IAFRe2dwLOhcYjdm0evQ+wn1opeteq
TSFTef8/Nq69hjfK/ii2f9VFVH/1Lfrj2GkBtRI669/1LQIpJkT+/kKU/CLPHYlk
yBnbm505WlklIrEP6Tt/ZG6YFGXqj7Y1JYpDv/rzZdlKr54IuU8tJsoKjXEpVu6Z
7Afqv9ZEnCaZ+bUhF9SPFKbZwJvyyRORWRJFvXPDn25weH+59J9XhauJcqOglQzu
bpQwTX9sfzuuMZOYWd/9XZSOUlRcCPfSB/RFevPLCbAr6mXyY3PTnEEZ0etFM5uG
6M8vUxfBY59iNfxhDkBl5gNIzHCwHGBwbIJma9S5yHWbr82LVlm8flspwMu6lw5K
wTSYoeP7NNzj+3pNQzHDXnfYeNvO1XoMuZWkWUqM5aXEq7UJRosse/jztGNyb3qG
k52D/IXqPMoBOyml/DNyptVd1O9C7wPfOn/bxl3I0m4JbLBqY637rkXwWzpIYVBW
55PCpg6iHHqdCKQZt8U5Wf6PD4QkAPNeF1/uuD793n0w4b5QXISjwvJoM/kFcqXZ
7jFLXwq/4L/m6n8xbTaUmXjwCvSl1jR3TC+RBXjQcyGAvZOuh+5XjvuLAfYrU5wQ
SCyzzKDOcfn+U+r8YwaXiyfUuYm0DJtJMYarsroeHOJ9qcVVyazibpjF3U/J+vZj
+6mceHyEs92yFNIcPVpKpBcupM7PfU+IAK0bueuu62qy51FAx2wX56jAXIKJpYqa
A0iadlpqE1fogfR5+TpbTIoGiGH7DtngtMFGxz+YIDZRmMPOrwDosYF/zc6GVQ/o
FtRBZ2UQ/n0AAd1elM88HrikStqhcl8/DaTVfG7VEgNhek4/qSWtoFeLbGBLu6Gv
COY84ogumcWETDQi9dsPULg8YQFRlwcMPOHk3qkf+TMpo5CpeJj+yrVVaqmJcWpJ
XuLVOzpFqlFlXSCJ4fNDbY4SuR50kZbtUHVPvS4g9SEgvtkplrGXZk7UI2Sz+DAE
JLOYVH7sApWK58HiIqim1fsTKWpHmhcQRQ3xzzlxepjA/JyC/iac8rl7X+0Bam07
LWUd5A2lzEO9LFw5o07AjeL1ZAwby0AQll5A8IQNw/VuXJkKmm3ZQqO0Q0xI2x6Z
T5GyoAejNGC0bufDZ++B9BaYGEr3LrSWb6EtkoHjamKxx0tyuXl2QM31yTYFoNZH
gTM8J/r/jF3zYBA7m6D4StCagQq4/+dRPLAfcKEEaHhd6NwDVm+yt5avxSMelYlC
BNpaWlxkIz5xDtkGKphAU4Pa+JnYB//x55kdPLuuvdZyme7IPOtQGI6jWtWVjKfJ
XY0t05oK0sX6ZbZt9XcosCZTE3qMpb3nLA6kidDAs9URtI5ZkyVwAc1kMsKVhtvs
H/mfpoItgXK0g86aNdsLcZ7QHtNlrSLmXeC6T2y+a1sq21unSxsgopV989jG8J5X
fa2WIxTsMvcf1aULLwF6+RtqrrJxaJovActNMIwmBE9vi7HkyYvWnXMcjIA/YhQl
Xrty848LeU+eG7UQ7OxQOyGahCdw2/rnvZG0OWM0n+KvflgEuvqXaxL1EyApgQpE
gEsdQMqwI3b4YIf9FaIhSK+qb7OkrQQMZG56rIMaJpvApP6B/bak5SE1D4UCQk2E
KaJBLZdBzf2zmBxvW9U/ij7cqnOE9DXo66SZjOP+WRqS9zDfK6SDc4k4tNNkgPQ1
FmkGoRF1YyeDgVZPGY6ZsinhLQGlnkq4DNbE306UM6amprYLkZFt1FdFO+gSlpu1
Q7t8nrbIQvW+M0w+/WGA7XQzYSZh32NIQkVgHB3jIT4O1mXE0vgMirhbKuEP43zm
KRBTIYcNu2Wuuq7N9k0k5nionfzrsTsm4CK4JzgaZnd/GS0G1/B3ObF0g35QQO4E
VVq8VoAAP5uMgc5L/SiLxpRzyO/rR2Z7yIQexZhySHDPiq98E81fwCMlJflxpovv
8+DS0+I6I/Lriwls9IZPR26oi93Vo1xZcRWiWK3fzipXfObPJJbfaZ8h9Q1LpxXn
TTIXgWJQEa9YZ7knSgxcRGvl+BCp1rSKkGjEsMmkOp2uLIwyp28CceLbXGT22+xR
iKpo1qZrDUEbSiVe10ldN3o/PlAZfAfzw5N6D0Mt6Kj2wqi2Dt3pxWg8069chngn
TTP12j5KAsYqG3hD08lNbf0HDfRRemhKkbl4Z3Pbg+Ip6eghWiqrH7BIzOQzLIDJ
Dk1pubNmNrUcM1NJp+ETy/u3f2BJSqcybwqyPkjJxu3XJnUdiCOi6oZ2khGuzikq
1JXxI8ZWefd9Bx+O++1u+5zDsXTGp5LRkYhOYeEbxm6r9LXFdZdOQQYWGYIpYNf5
Rd71Cf1MP6O7ATNJ0B/V9uXa5meWDwI0+5LJMduJeLQ+I3d2vIHsrJir6u10cJtl
ZGeGXwDcF+nEWVjTPNSU2LjDk7tO04/Cw1+nz4+Re2+Z19DfiAt4s1vRhccNu6uK
IpPZBbWbirQjRKlkIsortzHsyahJ0vPf0lrOXJFIoYVtVW2Y983aKnYYU1gbRzEj
mgmYYlB9ZBR4lysSBwyXrhdvWQNTkjufrk2KVfAhpX7ImLwOqdFmQwaHfcKwv8iX
2FLwomK2UdrnUEEie2GUalGowGQk9a++szlxxDUoYfKm1wG8Zg8CqHHm9iHHk8W1
wpQJh8YWSEMUcLeXkDVjF60qBz7aZKf/xHrq0bI6G0dxDamak4VSEpP82+dNtljv
9j6T3X9IlcAH/bviBq8idtduEuz9oN439N/jaGQCscK8KWLRgawSC1doHd+7VMij
/L7yvmmSus3pouYUEdqUrK8SigrvpcNPO2CgHXYCFhSliQhiAlAvB0rdYkThBwce
LTjOA+verRrhCk3yItF8FRHZ2vq2MG+PkZzPRPzfxuUVGNppMAeJbaBvFphRAesV
kFdqPF7DQfqHUrObixcLUXvv+dr9a+D/C+UVmKxK3s5oi+TaAhGnzei8vTJLA8Zu
k0ICbaO9f0M2Bf507dsN/q2WMOzuarO+h2NeM2t8itulikbrS9pHOQpDz/Z8gpBA
mmo0aOnYE4BY4Uad8RwIpbFPK6H39ujSmVep/2mPV80MgzZDlo+0s30CV7b1j3dA
rUIr9PVcAy58IU9J35vJ7VPVyxrwvjKEvudVmkgy1IdUpmnQdixQ6dyVO6P+bdlv
muqr7oL6zqGPWR0ataPkMhMIOA1Txw26oh0EMULcAFsMVhbWeGz3H8vmsvdWDu6j
jYouwp1iZhDEc9mLYqcZ+LdlNLvQguS+xYt1dW55P3AXt9/YqI7QLZTmLOq/t4bx
nn4YmGw5ILunJq7kq3PDpAIKz2ZNo1VBIvuBf9HyViWigQV34KXq9LflDUhNjH8U
V9rncX8CBGWSzE89jX59OkqLla7w+A0kf1E5diYNOM/sNv29uzCHn1btYBXD87oE
ER+YLw/jygTQVXcdGEnAShBToDDC6QQG0bQGRj7UlqkAMylVVzXoLa5FquLITQk1
yNZgtaOF8QPnxYmWbD5ifRKwh2Ou5gHZjbclTvGwuDfzUvcKVVFIT5ST3W6+fmNL
7FcmKT/j7SAjeNdkiwIuQOzROBzjz3qeppB0COxgKbuApNopenbER4r8Rb49Vzxy
X5gqmRTpO+rf2SkipJdGagXYdwjkFVemLfjlXqJJ7YJgjY+yEckOWPKNXQoy1XSA
odDQKNNk+x4D7uh8i0h4ppqs/E2ZESROc27NsLuH938PWEh4AVnq+2uoWu8hwH5R

//pragma protect end_data_block
//pragma protect digest_block
sibJFcswUoTDsuXNtDZ6CRFh0Hk=
//pragma protect end_digest_block
//pragma protect end_protected
