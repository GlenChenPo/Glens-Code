//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ioxRnEctqJ7RtGnXg6dh9jZB2QaKrTZom2ev1RugP74Fvo9egY4eeUxzWbq7E3WG
XwyUoZFyMMXHJKW24z5+FnfOd9SkLYysqae3PCsZn4aaBNazltR8LagN7P1inxyZ
PjsusC5R0uS0A5sKC2+ESgQWKTEVJzF7KvxzFSto4gvSFiKUCvz67w==
//pragma protect end_key_block
//pragma protect digest_block
INMyomAm3OYLXmeN2UOGxQ3tBGE=
//pragma protect end_digest_block
//pragma protect data_block
1ZUoO+E3i152MWnaS3BIZTQaTcsAUtp2TXjYjWPcP5ahBfN69yU6tpH9EIEk6NUV
tLxEIhD/gfMP5P0oB4c3SyEG7RGUWxFJllWrmcgKFgzNeboWIPcg5kyqR8c5SlvM
gheZJ4jC1vLAF+vGCPvMkalw9GWjHXeiUH5l0lvPPRRRLSsriod4VcoTs3ym7aw1
rlu0/fItchnfDNF4gF00Z4sFc+NNZ1zPadfhsObcD47XNNTju2vzKfHrULrmcq4U
FVETPpktw5O5LlojzrxIhl6b5CURULc5+UZ5oqZfyKlwhiDnu7O4DDCX0/mYaIvf
QWDaOQhLwtVzt5DOUhGkKg==
//pragma protect end_data_block
//pragma protect digest_block
RgBRXLq7CL5NyZAKsSJzF6S6Z+w=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
eKaO/mxoNPpo1QHAmkrAkpVG6sV6cp7xuFiNTWC9Tu9Bse/HysXQnFH9Z3DFRY19
ryqGWGHZWyFqKbBJNXN4mG1Mzcxfo1eVFoJ0p5RckiU190yz4R7GhSuZsqLdqPhf
zVwaDNbv8TMx7bsNDPt/GAJ2Rri01WWOMdvy1eyqkF9S/hehyG5YlQ==
//pragma protect end_key_block
//pragma protect digest_block
0/C1f43boesIeFkYwprxGpnSK14=
//pragma protect end_digest_block
//pragma protect data_block
k9VGVcOfhDRT4Vtw5pScskU2cEatyQjNRXJ8pqXpQ6iKr2URtGXayRAhx+tb8hav
8Dp5IS0LlpuZDfeiCcRjT64yV0ZEa7gZ812Ojysvk+o8Y1UZLWmvD4s/gjnv1dTv
69lZPWQbLZLaIDfMXEWa53rZGNIFfkxpv26oDJcVGimk2ywWdCHU5m+FD87s0flI
gGMrCj3+TVNfs3HWZri2fYV8eOrmAunOtBBXeV8GIUTiRg4kcuv7zEJu8AAq7fvw
dDPptC/wFgiS9vrzsz855cdafnVklDU2XUXTdjPeDGNMzwUdR3yKAty3jFiQfP+K
ZvR5Zwqwji8Is9fTgfS71Q==
//pragma protect end_data_block
//pragma protect digest_block
G6WZVCoZ5y7131USIftYVnicZ8o=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KMV8KX3Z+Da1k0z7o6VkaKE3CH+yPd7xtFMZHDT1EC3gHxIdW2MFVWtKZr8BDu/5
uLsNrECjAyyiVqjlbgmkG5BW65I/TZmZtevXju/3beBPb4lS91hnpVp6zSJThMFQ
TT5o+7oXJLjKyzk1ynmEv0ugSEGltajfFYM9ns8Y/tHjepUlRlZxhg==
//pragma protect end_key_block
//pragma protect digest_block
2dRkIrXBafjueldfyOkYFaNfyb0=
//pragma protect end_digest_block
//pragma protect data_block
yzcP2poYaBtDMD1AVzfunuzJWW4aJYumMckTZ00PZUhIAgjzw3nkwzJBUPWGjMv2
Bqii9/4GDYQ44NOneqPR+wr1qzesX44RfeDF972mXKzsLJRqYbDwy3UiGbjMgF/g
XIUqMES8QhHJq0CcuukBKInkpIpajdo3nWk6cKrjqX2+QcmOwYcUfEqNz3gfLeM6
0SYRVstPU+hR8PxwBhCa8/VQTSLo8j8aBYDzbHD3IbEH810pF+O22cnG/E3D5F7X
S+AZyYwQOx1IT/nEhtSTxcLDIoWPv/5GF8sa5TBJgltjybkwjGyv6Kbfnkmkc9Fn
M45aHmQ7+A2Z83aBi+ZR/DDh/GbGXE9ZMIHwq7iquIzRvOj+rTkG1Om2RArB5o2l
FPhlYdourRw/f9dJJrmouboTZiS8O4cKpGWA4wESZzdJr/t1AB2QtaRV+nArlQ7j
shKZ03CFcPnduoHdkzFevIWSpAeV3vHNQ4bH2alb5nmgxYGKs0456KD0pk/YYHHD
O02HMElV66iV4X6v4goxnZHcDB8mjeJsCZmsch743FfRDvM2Bxa7rln2P+Jb5sN5
IElM0vOn9Gdwb4TfawleciwhNW0eNhXsa1vUWeAozuJJw4oDqZ54sxRDfgS+UiTJ
3axBaa4aQvadbsTOX38OWeXu8QjCOzOxOpvZ5uOy9hjxiepuDjsoHgMPvFCRC79X
YKq7MHYYGuyZYkBnepeKRQ7bYZBs8AIQD9yc0u6IY1d9bl0lU9K+N0qgWQtX1n3Q
DLcoqQGym0Tt38XLAfu3iAGPLZuRPZ+ASE1sEAelg0WEK43/4Wg87i3Dp1ynGNSs
mBUnI7+OQMxhwp32XZdjr60nxj4qTk1JpHs8wReT7htPVkRDo4xgnd69of+wFNwa
y8n1/9Ja9NfzdrEpF8BFa3d93NDjWewSlbSEUUQrPpVqmZRNtyquZDwue+qacWBP
Wk9j7v5sa6zso/fkD+rGyHLktduuPoKgBuIIZ4jfMod/VdrlOxiSnyXey++K7wd9
mBWG7UAfDYvpf4ydd+Lxlgwnstm0SrL9rRq+ziFd9DNPeUcyKk2UeqYR8vqSJEDy
o1c0KJigVVhw52nufybv0sKTe8HF1M17Yi38xx5o8+8dwtkiSiwr4wDRsxBvD2VL
YxLpUDPwMnXC2lG3Qad85W6LnXWLFfInoD8n9H/NrR+laFSg/EuHD4XhXLKknLQU
LH4iRR93boL6KKf1RAATj/7PHKrITCPNL1k36NoCMoHnjNZCr2yJJECOlEmiBxGT
VN0je0QXVm1X2V+byahrPB031qbJ4B+VeMFZLGpDwYNiT+xYKzbuagZK8xWGwU2L
OJyLgS68PNyTdI0xADpmlUzQlmK4u9ybicW32sj3HaD3n06r+5YLCd5vccYY4Usy
s9hFnJ/1ui2EsEWQgtdoyQMhst4OLrbov7xvhdwKaCJOfEHLhSmBEGSY63kJW3mR
fmCFcs+sSZ+ZKwMwCGDGd3pOkLxYTMq0Yiy21vDTGWJhTxadXo5MbpwDT2Ik/eDh
HFxVor00SxTkbwl71BdBIBXCmCEUVKAlCpgk3fHIjkScGHp3yO5SRlqzIcjaPte6
8xM56YDqFmkTysTPHXBUHeWgeFKVaH+5i7J3ErdKFQT2M7H1Pu2ePCEbCRqTU8Xn
l5jw+cwPVTKGicoLNSTKgo0kpEVa598Cep5PybNsVdGq7fVrdkW6DWIOuY7nAQqn
3eYpymD8yJjhFy4fWxZa0sUsOkA9ovV4rh9jCYyjLxF0jrinukPmTQYtjmWr8Ywn
ndIADbLz5iSv7/r0MdU69HeJfACr8X58SMebD2EE1dCQQZsJUKP4EIVbzgl8B3Cj
r7PBMOcFg4T+qvhUwyJDt1qiMVviXHS2FY7ldsw1h8j1IgYGO8KFs1I9TJpzVNto
0OPERIhEg3zRhDchvk6z1uDhCum0oRNEogKwEI1exyUMEwz1L0MgULjv/ooLC2k+
g11jMh1Tbv8V67XvVhzhAs/vuk7cZ7U+Gu7lXMZn9000ENxE5u+lkw342Dx5uVOO
7u2cVX8+7VN4WXDJDJCNchhMBtTNqI1rdh1rhmg8huf9T+qPOF0Tc0MtMACyJWTi
uLwaPUtzBURj55/eG2m1P9/5KH3YEGUuhSE8SmK1dMNAoKGYV5bnu9HY0lpIiGVm
sOZeOstoiOA0fEFLoIPAfUXncefA3mW5qycFh6e42vFwk5ZoTUk64p0dIutNk+kZ
97v1goX55qOzox+uI3xY1VPxc9q8+QLepGNTCeXlRO5jYZ+nMza85+ZFxIBIgKay
Huf+/Zg2WifAkBeMkts5dFH90CkNNJuQg+RbA9UKD9Zp5npn/LoEL05vBxgDKAcl
TG++lhIhBLDC0L75lnSDCDPKSEylbhP9jKdD/Xls6IE8K0URlIcKsR3CFlfy22FE
0yjmfxhDl7Ulz4JkxEfItWBxSbQZXgGq7tRPYPchYuSEXhKusdTetrUetL0otI/R
/1HdkPQ7ChHqX9+e0nDxqc7kyma72j3LQbTU2KYw0FlgSfNqZWr6U3dtSbgu1cBn
2bMvon552LnSwFs32lFr6hDnH+ISlFTRgi71nn/PoDG6CuFrVOv7XtrZyA+1bzVT
sIW4xXLwUIECrEzkKZST6U2yK95w1kWJXxxGxQH6X89berf8S7h2Jd/GWej08ail
memmSExnF1oVm5FQKm0svpRHZ0dHeje47CD6O5Nu7XD8SlqIBssQKHh4G1czsV1a
ksABqAzhIkA+gwpA6pYZi3UtW4M2MD8qlvL252ho9sN62yAlmjJ7UZ3q0LRQ5A0L
bIoqdUjYTO8vyKiXZwUbcdeKmHGiKoAZ6L8fCBxGc23kBqLospCeO7TTXmzWzyZr
NOgPrO76do54r0ZyGVoerVD0cUr0i4RFaHp4ARDvWJi3I7nCykO7DFeYozKB8sP1
qjTqbZZgPZhnNbeUx2iLLKuDhBoa3DkcavruV+dV64CG24K8mtLTao1Y3+tZds4J
UBt6UfNCeMXrwrnCgQeUkht4/EIrv/SQG3x+Jv8FEt8c0rBlDvY3frSEc6pAstlN
8JsTuQ5ZSN3i4ENuvvWPqMwru//QX/chXs5ExV74Hy8XjWZi9eYUMdGRxcOgQHC1
4ZP6mp8hqIXVjsJcsMi5IKtVKExzpySMBYlQML4tTFF8u8Vq+bcJjnoV7zTCT0eL
aufi/TItszS+Ra7CERFgGSbELYBBib2CxrVFTEzWyhWPSkkDlwQh60a78fnRdIuR
1Tqri7AvFCueD6tSALJfH09LPzyams56hIpdsfm59CSepUhOv4fwo3DiaMMt9X54
fdbrIlTO/vGKzoSAflhEZREL93WGWPD1P1kNO/BYEiARIAPWvBAAznljserBxvdE
djzIu81PE9tKpGXYDE0t3xsa646M5XT9XmGpPpKmxIray/yIAaG7K/d8Pru4FbsF
AVcDsF7zXeasxBGHrnsGZBDVmQmr4nOlDpn12yQiDGsc0yLLiznxGTqg6T2kp+Gg
fe9wNY8EVvRci1KoF70wxWFJLrShELegBv2n5zcBoGUieKEi8mzKLJgJ/a9V9QSt
74NRHu7qjQMHmU0YZG5JFlJbRdP7atCudWzMZRm7z3Uh+Mby1NkUv0++FSmVPVFe
PrVpZ4slvUE7Aa0Ipig2n0LVrh1RU0mzlW+84VeBRiHwAhvzxeQO3fEZaKj5kJxy
D1hEwCA1A8ESdAZQISiCahMZObyQsQBlTp3kRgrW2eRNaOo6kQjuXV9eSjNsTQi7
yeiA8tN4J8UQcS3tI/CRMCWnVdOAD+N7YjFd86vetjGaieSbyZMY+oehDdyTjnZf
G4+R9PRdp5xsE801ywUMHv0H8lfVkP65nnolJPHb8/n38UrAboX1txL1J9CbvbVT
2n2acHt7nlDs82WwZfha/wyDNzYCNeLJtHvwB7sXbSNaBBwc8fwtJTx+pV2kPmWH
WdsmP0qSPZu582CiHNmCW/v+vwYO4/N5mmQ6CXSgbnkObq2Wf4UbyDhmJ5GzYnMa
jGWihzZILEShiIfP2jGBEPSbfZcuyJ4AAeUASuXb7BVg/lrj9J+FqZqTOcMhkC/v
c1kvNrvIUy7vwD9QlpgSHcO0BCCX9xB88UAnY0TJlP42cZ2DMkslMCc+YzSourVC
QMR2t+a/ODv87iHBDprxBqa84EcpLY9p3ZsgsbIL5qu9Sno9xebZmt9tMxQQKfBj
7gBf+GLs6aIhPQMN9+98Vkap6cBGfUOouOTnRMgc1HyQFES8IYpGR2gODigvUX5Q
oiKB3xGiFlYIDJ+a0FZNdmP0Q2Rd7Nq8c3Sl4X66YVr2OBFuESNcoeSjTrHylccr
HNzFX0eZRR0ey9GZabAoHzNlar37FET4wQmofOliw1opFkUpQDuZ+r+o+S/+RYCa
SGoMWPMK7PItrn4w2diRkXnd3qlK6gLkSrPEG+JOBswbiq0HrvfePo0M8J2KkVuO
negteqrIBS1cbfuWl16ljBwXEmkce2r8wTi1P9fMiY/6ZPVM679YeQ9++ubLFBbb
pcpKhf3F+J/gUtUsKqffHhr5oC6Y4Fa0rWFwdorhFZx92WUwwnV6wMQ4eYg5Y1cK
COU5zTMLzJHTCIWbBQ18rt07rd58Kwqzpqk/Ae4C0eAFRwIQR9bg43XqF+NBVJu7
rPeKKxKecKZSu+xtpy8bznZn6GQr/IDMjCcUcwXlRVLMFuXvRveovM3vO6SPdAlo
xRIy6h1/qP6UeLedRIeoWeEi4ALzsl+Ce0rxh5g1UWIHrlzFAHiP7HRm7zhy4C/S
8MlYFEhXrMlPlISZaYPjuvyxkyBKoC1aHLTkMNUdRYvy8LoAF7lRaAQJcVPtDBJm
62HiPg5eIW/MQ9NwuZjvN5tT40QHx/wWrv/fCrpeZQxd2hIwYqyi5awfZPrSklZZ
RdBYzHZx1/WDa2Sy+ay8Q3oVcHniZC8cLWnqm5ebSjigalATcUGH6PKDMGhoOQLO
0TY7Gkv1sgmDyvO0aql15Ao/PrneF1x40quotA0LbZj6Zeq9KYojjRX4pFcPAdca
vCHMTzN4PcCcUVjR8m8OV4DogL5rCB5Y1dtP7GS0tN7GcCH1XtIzt3vey/a+ksvH
TQosCW61oms5+BqCQcYWHzNcBOitaZ3sRCLxiOQLPZxxCNSVMAaCoqnLw69+0VdL
aXr0pXvtaciKTLR68dVLa8k/Ei+OIQOAGdnNkxXzySQARwZ9u+8CGWJzNwVCzy3p
hKDH4NAgflvMfUdE0t6vAWgUSenlmxkbW3qQfhxft34CierS8525E+4YU57yJKMa
/5biHC7uIjGqgmA0l1Zf9pvO3PBlqclUYAnnKgReiZ3hesXsBgjWZTi74hU6VRq/
rcZNVrnGymqPiTsTLHAv0PqI55/bva9Lk7obaCqcqjbgwy4OW09is9I8Y8QPx85h
D/sA6RayDc8RTY762G4R9R2F0wKFKgxMl7deocD4QOO7epw3946ECqt4z5FPOA2h
Gs20Rh9Fj7ONUuBm3vI7zwh9E6D9uHul5ABlXS7guafUU9mkZJ+pQK9nxtBQeM6O
IlikJ8dkgRKMJdtwX+fDkanXfRHg3pSTcBasZBamXY9iePqmHMziL4ILyQDsUi8s
wcCsaMdEsaLztW6BWV7FUK8tPOFCCVmHPT6BH400El1Fd3qSf4pM1wg/nkBwg6B3
cAVCeUZLZ8XkVOhxewrgV6LQHOSCpf3qwoDErh1In8fpJ/V1YkB1WGSzyKDZkiQ7
CuYzOmqAe8YoevCf0u6Z4ZIe2canjQR62Nr3YMKSWCInDLI0evb8yX1VErHPc/4T
XesBihY53XEvTIpbKnn55qFAewkIFXe7saIQx1n8/vIN8pTDcjHRQeOLkf0s42HR
bnuxTZ4WiAY76eRp2D2vmWg+CsGTHbQQwf0yKJQoU7z/d86A1/PzzrlgBRJuZkSA
nhEnIuYJ7BXFxfdUFWjJUrz9qa0eMREvX8etidizA6st6rSO78UNnKJV0teqmzwp
U3hqJlMan6bcEt4I+KvpzKXdG7B/TPCVB9ElgIxURxkZaBCup74G9OTg+coMHX2K
H1VdtJr6Qc0W4mumWd0FuQK4LEGxiovXiS3Qw3LcCU4jQZjdf+PwRhqdklvPu5Gc
m7AQ6FASjAjGDsfJomvsM6SQ9szIsuCh0s4mWnJDRVU69fmbQ4H/Y07y5KGnwI4T
MnIa+H8whI/qpKPMvzET/V2bvL+/bJNQ+ERnZXFLHvrkNGguVVUQ81Fp5uG7nkcm
A4oDacDrQ+YIO6uSXBf2mhNxk3qwy+n+SXsh/MSZb4jTaSyX/d8zqkOj0ak+FnpG
0tTVnNPbSDJMxgWUWoP0vMyhqi7zSxnEzH3iGJs3FkjY8QPmhIBZUp6DcofkIG3k
iPCnwILFpBt5P7Ga0xzoYDGRojBTnPIkY1vaox7Bc7cflGPlx7BMZ6pEuQZMxqjI
FrQK2wA6LFHMqesrGIbc48F3fHK97g1ACTGrae/Crp1Phf+kG8hqfG/4hRNtoFdD
uC+L6loySJYeyqjcy1dCe2voXcmm4upfAit3QdfEJWwAuT1ppBXmXKLFS2Vz0bkw
rM7IpXIIzzorcgBQLNqN0L74bPEZkIFFqPvq0sfqFJ3umQfP4NtlupUlorDMJZyI
fjk9ft29gHUYctBEzECxl4je4SdL3dFnYIdbi7WYhiEbxaEUlQt28cMcPvkzzt5u
NUf0UNLk+Wfb6a5RH1s1phuJ2/Dckw/AMJZ8ndaOYmJOk1ZyB8e1ql6Akbsr2Ta8
ASJbQyHwqnfz+Faz9bMrP7YeS8Nv0S7rwi5VwOkYlTIp07f5yXx6J/XPtNwNCSck
StdIjUTHiiaq6mjYsFHVcPtvLVwA21aEjel+vqIrFeXPiB9bYH61AygDg4PclnI7
LomyVLmrOwHEem6CsgYE9FyjSRp8tmB/gBO26iwt/Fzn1p3xR+NXuZXU/ZLE4y+O
BboDxZzZNTQuPyhT/mWYumhLgE8+DvLODcconsgPsbpLPHXK7o8gnM5L/6LgBMJX
PK/5t04POYJRXqw2waWwHL9dooDOYLB9P7I+CrlSfy/AK7ilHI/55mJw5RfxRi/6
qSEGHOQGCXYjHiM2JcicbB7IbVC4JIG2jJo4S1lcADMFrEqsDW0b5P9mwjJNRWxx
pv6JgkzdemXmGh24ZsyK3M4mfvhnYBZOmy+VTjfs9fXf6j/eryQOYc14zToVBXn8
08EqDb2PjmcU1zNE/0xpg0IgbRFjLnqgBghrGJZ0+TPjm3vY/JgzPgupUn2n46zu
NwpI622bQeQHhJozLj+Ppo6IDTCVb6/9H64u0bLSrcURKxbE9rWFQiyLZgWdXcNK
IWyBcT23Xcz4kX8pNUmmX+SoSce773f6f/Bgj4fqpEdsHvuOMLYLaZQkN4XjBthj
GXro6giey0IPybnX+EFhdD1/aWaSX5mhAy1LxHW5NsQPn5lTYdtqryGGv2gr2P0k
74JiMeZLaPgumRWp/dtLvmEiri7tKIKFs6GDphYAj6REQD8a3rZALUcTKy6dz9ho
IIFIKEWKLvJNqHMShj530QxP3dYYlBIt2Srd8zfN0+XWyTvSO72q+HrWv4cn2KDs
7EXhGe8Ff9ElfcBL88kB7K1D1chrLIVKvIbA72HT3cFrKGsFoVNebbDLkj4pKI0T
KEUpdKJtkXbwsI7962KLIn3uajPzsGu6AX0luh7zZv5PeeVuebvAZAFitBap4JVY
X2bXJpG3WFXOnLwSVVabKz5FkcjsuaWLNNTe4pM3RLHOci0bwcUFy5+IffQht6CH
LhJw23sGXDd9bm2hNRO7Dzx4CNywYjAR5WisMbRgwD8yYzEbo+0Rwnk8TxRwHiy/
LWaRDJxpd/WRfIib7R2Rh28zcLCNl8zQO8/z+2Mr9GtFgJH+X/Gbq4dnW4YMUif/
1GTNaNiIj6AlCRCk2Uq0Et3eRfC96N8Rt4VUqzcw0DotRYZB9NwJlXv9UrhLDi5G
tp5iK+z21MXVAdnLvyccKNYyqIvr7uqt1XjdbBy/lHaAF7VFvU5bbSddyh9oo/hG
0jGnxjIuXJ33TPZdVGVR5xDjGHp6hQj9PJ8bLEIJag6dfdKaPMVsB2IPJrdPmTFX
IYea1sc++PqGxKAM4wOay2FZknftCMtfePoUORP66uOpm6ViB+CfLLYiHM/siUuH
3/1suRSIDZbKk04cdt6cJcI0zy61OyLo419QFh1IuPTihiPRb3Lt97OmDmb2FwHP
Cer+dpnlOA8OYJIPGrz2ura7IhvQU6IbYf9u1S8oQk8eCDjd9jrYK7dHPrUb8FIq
oYgK/t/T0A8dhshiMmVv+iwVvauv6U5vQ3jhuT4WH08hAyaWZ2qbMGRs0YEYwj6Y
GHrhe2C1KINJS+VlSlE3/8fzmdRBuZBkIWFIXMIG3ys+2FEgwTX95F7cTz0+WRbm
jd0JwpZuVH7B2t3ns5OIUGN60gW5HMAsoPSbtUL2UYo6aRM5WQjwilWThE2C7XrK
lcDBseTePxRFEqqghuhuepAbqUtMuyr+kNPihIs8uRo55p6uzPEIhXS14ff+DOky
/aJvqfNLJpPOTG70mZZMVK7ABzZctWFKtj+kWeeKBHvUsLxCkAAxyrNyCo8FItdX
viBfNTTJ0SwARziy8T3xmNx7sOYay1FkUATRJHF3YHyReZj2KnlYXv8WoLASrUhf
c2ZAbCDiDI8WmDUjXZIQZmO6CHzCVNRnKHo1ad0/6R0+tQaJQrn/wi04S7wWNdgJ
CNvRz0QtcfFXe2OtN4W8XGR8+6xOfV/TB0UseC37ascU9Ve+ukKz0QyWmuLOOdFd
xeDZBkCw6u8BKKtm5M5BSaCshBegHob7d25pxpP3PSVSNZCyl1gFSU03ax1ZLokC
m7ZEJb8SuqAt8MhCpW48t0l0gV/JRhRtgJFwdJI82QKP6VNLf8h/sJwqsJekZCOb
Q7YNEpFGazHMPTaHkcG/KmkgFjthGSrBgOj0nLRepIe+28rYMjwztih3J5Kwx5Wn
o1gx6NSHQomfhp2J8VGE6W3zy71HeUVE+qRAbAQJgbfuCVThH7qDS3lZt7dpFuzB
YPrl1OPBtg7RBVD0PqVN1C26R81oFqr1Tue8ZEvPv5+h94SsKdS0wRnkk6Dc/vp6
51Y/elbkOU8ogU8HecIAN240n5wsu6F5ifTaXny9Ee66buDeQ5qFgnsbVnYmsfQt
QqzgnV6UGV3pqAU1z+Op3XQUcG6ByKzOMjpAYf1gfEaxLGJQfr3RxazOZw7+QYzi
oN9ADda5P2Lz58EHW/WLChwOjvaIw316KkzLhrGSZRxFGX5jN1B6OnvX9V2pwyPp
SktQegOrNyHgAx1OXtLLJp6pBHfTM2nYPeblF8+ym707rrFPFipB8mvgOu1c8Dbp
Gnwv+KqEZaZxYZa2xaD2ZL2eAngjT2t3Vk2toLgNhRx9Zc+AHHfZChHf6d9jA2zb
dM+eb/sWD6MlPSxVIHPra6jfurM14qOK3Kqc5iwWvFFZSwQc+LU2UtvwsTEToPIu
hiOw7PzOvVScnKDu1IzHYkS5SWGh5Yakj/v35WEFjdzvgeajrmm2JNEdfK0GKBd0
yOP7FWqMHgdL+OgYTRldc1jUkur9wz2w5cKJNSOJNuEq28b342N0GODJllSBGMbP
oiyclP+4/zUubsis5Idq024sqDkkbrp7q59btAIf1K6IVVQDU1kYZ49yRnWRoxGd
WS5CJrF6ww8DLsWv9hf5HeJzobFyhVBUulCVGIHk84mL7b1zNf5EN5EcuTR5mFvH
cP/iK9Fe3PJ4zwxbmJZ+/HrjR3ndkHebMrv//nOAipw7gtPNg5/KLJ5fXqc3FrSc
sFIsLiP6LAsnJnccWQXb9CPlzah25ZNXKEvZkffMfPeD7/q8fteg8T3nU8fSSLO7
eH6qAfJ60EcFdZTKL3ZYNhLIm0dMk8hm3PRrrdOrNTxmrjtv83C2B/LXu23vPg5Q
hjIGQabeYD1eH5wzEi6wF7R8fFV8Fx+UrRkpYCCO9M/ibUs+FcdylxsB5e7h0LOf
0ENwjIWSdyMlm2cYP7MoHtwJcrhjZjF0Gd54+OPmG16/uI4cq8qdyFJ6/aUgTrcd
0jlxQNW/daIJMa+v4UM+bEr/rua8AxpyVODJbtXTr/UupN8QNhZ5bpL/FEeaCgno
Tzj39eH9tfJJdr27cBijbkUkVQUgMz2Ovb8V6CUKeEv/5JfHQBaG8QoQwloM8gan
UL/3O7FKKhivt+D1aksJVo3zWC9l6GKkNMemFbKfv/Yyx+CeXjuzWtn1dl6UchTF
fCqKHUzk9ekispqwWa7M+EUaexpxGrACA5vn5oGrByffIJ3xCp8C+OwoZ/FMHEz+
DZc3RyAXNzcM3M62VPN7lJhEFKTqZ88c7KnSjHc6+4cHZYTqHGTyNd9rz54ifwPp
/77IPjoSqH4CmP15zzSqp989YTrAz0WyNvDnlXDjTDiPFU0f6qbNm1AnSjCD/OjA
r6fytg9LoU4udvXSGtd/YBe/lfYz+wY/UTJxi0ylJ/ODxE4RD9gziZ/49jsnNvyM
5tR/BOz7T0JRtPZAmzykFQeFwEocF7tj8iurXV22QAK1znTRV5NuzLGsSw0Lm+o4
HfqBxQD9Q49gLqmmWknGqUpteIXdlD2Py39Ngd8PS2e0D4vErisIaWLDdn3LEwl/
ka86xot2AZsXsk2FtREJlTU5gugdtvhI9r5jxCPrBuHX7R4VvnB9VIlKhnBeTfxY
orDX+nLgKfnUgMWD+SCezonOO1qqYTt4oIs/3XkegE/UQe77YgU8FYDjoudtb8Vr
ZTks/3qEP9wJtrs7OE6W8gumQOGSTxMr5AxI2TJEyhz3t+BLE/XghTtJIcubvURr
TVSYYHJOcp3MXRa8eD/DbNmRG3eP7FIxSveizjho+/2aYfFbBFuKqWS+I/HYG+88
17DpAj42DGKiI46G10g19eY9ecyKgTFrt/J2tNKLr/Nc4tGzRP5lRmhZLRDZP91Y
gdrWT1TDzbKcyhfqhjjHId3dMVdDTIBxmZF+PrTqR+R1UOOb0RRY9q6SBavt7blb
OiXOX9pr9xp6/1RG1bWRu4ou8eRI4mq0PwJ0BCC5FkPrGkZAImVUDB/atJqWGS7E
MVUivnNjzb0Klg506PAdzM1N86Gab/roRtS+M+m3/RYJR7pnhYeqTBCdAp7pqGj3
2M1nf6/YGe2PukD+Kxgqz5abOvcvjoZcC9MPqQNzdt09GWJz7Z03Aj69dg0EGYou
mc+2Om4jU6+uvpm7gs7zkKUOB/DwmnE5aDNzsTijyxZ29tAVH8fxrGaFA9ULcoWc
6XAy/gyXGRHcGBU6uDE52Am0kc+Vsv2sk5ihNlNS0WF7AKegFjO1BNy50SPbNtIV
kjhfLnNDtEzZV1eaqKPWtj1SXDJBcMdJSwOtlvppi8AMoDsCbf6JvZkJvDtRSeqJ
N7TdGZ+RUxorsyiDQYh57mGLL9j2iVhZ8vCdgP8ozsgdGTP7wi8thPpCLcVDN+ds
oMLMDmTp2VuPHlDacXMw2V4oPN3GvelTf3XK3D/1BzhXoEMebY266LFC8SHD5mwl
R0rhi+IvMtkxNJo9hyyiWuggoB0WDhC8HuF/f6LL1Y0/uJHnC2sP9/dKl3nCBTua
LJsslNEyRRVzMcExf587FdE1OMOC9I6lunkFjyfoRIjphyPPaMmsgq10Y/ZE50W0
YB24l7NjcQ0kfm32tgY2m52zBE+CtKCHxDtpl5m3+7tdOZReXrlX/CkOgQ2S2T2H
MwidLGRYj1r5QWvaS/jjJChTvvqPuslca7Sq7UHbdhsvkuzSYzI+HMyLAoJH8gre
8dG+z1BHsuPrpxIV8YRHC7s/ZF66MttICHnxP9EqBsOLT+UOoRniq0nfX7Sx/5Ay
jccqcKssOElgyweKxcGiv70OFkun/Tzvd49QaB3UcnohuXGb2nxdAFx+BPl8R5Ii
4YFL6xQprkd0t2b4XOouU1Qrfv2PzAPoRg9mSrf/wbSoaX8dE58ji63jxcKoKEmj
3B9rYauZF+vWgUUllJC0o4fj2F+dZcpw5wL4HNWkYLosAWI32ew8gTHUvpZT3jXT
Nujanw9lygE0XkAxYvalMLbuqPdvqh7tWCu3RBXwkHqAnPoDg9c0H4zyDkqy0isW
U5vCXapH/zWjDv21YCJNPWlOUwfyB/ctV1dv0xRYpeTAbMtos3MyFfAhu+qMeRvx
gLQj2kKua+aXSHkv8y7NuNPwGuiYRkrXark5xFmzC+N4SUgQ4iGVYTRsRWWDZi5e
9Qp2XpdhHwJzWAo4YYTMIwo3lQRe9FMklFMrqg2fAHVkEvECzgZnz/2WoxLWwMBl
UbJqDBh2+0Y3andcg1nRHk+iE/2OPPyujthBbd4fah/Vf26rAA1UKhar0+5jOWEb
MklMaXRn7zuVNvOoJrmhCAL+noh17Cyj18moqCTjh2NPKTdZdNlwBuddZN6n9I4A
B1gf8h14sLQ4t1eSz2lHTFM+UxbTrVHvmPnsgOEsRDYFon+3iim+tt7fcFIidLRG
pwBowr6Odhk/5BdTEUpv+JhWagVyYbQuvbIveO/voLaTCjRvVuzwWo40FbB2E5jg
N+YChzHcT/Huekm058xpoaAGK1tp7whwOXphCLvyi5wIE6nwX8lvnV8G19P01iLN
tqRATVAQu0vuRhL4L1YKje2hfKOnkB3mvy6bku+50ECTzeXd0dtrViaDZOAcoSKv
jjLZaADx4HUbk4Oanh/umQZYjBheMvBdE6xwcvXBQ4Do2eelt5FP2V3Ttt8Gruvn
DpMVLGgnxCsxyAzPxp9DgTMHmvjAaqInOFJ9AsteiWm9KoxxNyrVkr3Imbt1DPK7
rBZtP2e/vqPaMvIoXKa9pqtWHmOa8PxMkSL+coyWBJYhKpFx93/YmInYrxf1gis1
6CKCZeraRhUGzfAF6Pi8RS6ZCLiQlHI8GAZ8Uh3XDJgnXQvPe831cykT6/7oyXqo
NfVHZJaFfi2Qjh6zwqBrgCQ8d1e/AI/DavHlqOkSPcC1egln/4Dl7EG/YmdpupCF
XYBE9PB3//nkFLLkVqW0dYIQhr7I4PWTF2eQw0BqKylL1HDVUv76PW5rQc2e2hdm
eYMmU4y7dVrqgTYMf9LjqWPKVNdcQyeDyGE2S1rTS3ngoiUAm+1kOInqFWIyt1yk
jX6Jgife9kOZhI+wkkSfMwMpxskhsZKFzt+ypYPjWJRlD1nYyeiEQh++ziME5v23
y+jNCwG++fJbTH2K8fu2dhHCVs1VHH3OjZUWRuUNX3W3gAQ4HbI9B7vkQYmLe1s4
4MMvi23e3ALBqtfX/GVVCffBto8zygkE+nswe/MTkSAtf+tGFm9Cpto4vchTiHB0
J9vjvANTDPD7xvNQYC52S3urcz+xqlwnUk8k4LPKeONeiffJ5GULPP5iFyt4BNx1
4oJUNAXjcrpqP9qA2FKWGg8s/i9oxNcMwqmG9FL/XSzPqZ89uPshBYnopN+PkE5o
fpnAIyQL0EiIU5BREm4fMP5ggjhUG36q868b9wNvn7s/z48WOGy6RlNJ2L5Ykn3S
UaIk6mEQRJqdvMo+5CwXKl3d9vjPRvT9PLRZEOJGWYK+un0OoJ5kvNy84o2jrkZA
fhd59479JW+sq24tzZURtcexdz9YYVSUYfkMbEkl33miO01fu3ZvIKjj99pkPVw9
TKWTDzXk2j6LYu1FDHHNHaS5LJNwmnK7nJYsGztC6vDcq5X1y+aeBlqfXeXaA+cl
YW9wyjmDwb+Hh6pb/od+yB0wiEm0gPdgxwZcRXcXMzCZ3pK438oK6IDxQt7Th9QF
gpIgRROjpFlt300O07suw4GKPjCOwI1HUiy/du7+3FH2uRw7T0g9BA3fUaCuGABo
8BppSKWQgS0gG2OxeffyH0jeodk6MJezt/jRp6+mpBCklZrxGDx/JHDIUlJpEqo2
lQOKE+ZWmr2/gLXCxQXPDzBScE95i1fmZ9VDMZWMu0/OeyoW7ryJzk6Z5I4gEM0f
1cOu3nADgwx/D+zuqedCppYon7AtWsKmkb+WRH+2tIdW443pnabcfYdLFSbEM8KP
+erDzcBFfZbUv6GFnuOVtu+FeBH8b7aASBBecpIkS/UGh6D7X7kmURCQbxW7BHdv
v5I3qUhSqcB0lVVBkxehWi+t9wlUKWf4IkWUzwj0Pg3YwRufix8+ydv9vcCvEYI2
6iEvxhEUSvOAmNmqia6PFFpvIO8WrnXPRCJ/SDCCmcgYfmId/BQGCNX2lLi5dCag
hUK+CJ/7C2Jz3y9kbIoOwvguCpDMj3TkGZgiRoj11Yl238h5PWiFlXnuRlG5mEy9
P2k6jNsXrEOQAg9cqfdv6exU9CEHR1uKZD8p2VmIrJNCPNWF7TQiN3xIweiFWlDs
r3/gkVbTAM/G6WZLXvYEaRTBGr36XKZLSzZCmdcGpbaQNc+5ZtTDWVh+ohuAjpYi
2tuI6WzFH/GSFqMq+s8ECT9MJyZBY3DrS8bn2xqPFpZzNcwlEFC5xxPWOnqdyCSl
UYjXuywTIeQz4bgJiyFgBn//osDt0IZ9ndHLBiqtoBQiz56C5/Sf1GwQgGKP5jc8
+7JIHZQ2i5cUKzikXT8Iz4Nt+4i2y5x5JJyXg57WZoxRiAVchSiclGpmKWRvkR9L
jys1VlHUcgAk+jqL2j0CFoe2Zfd/CXh6W2D8BZPp+iCMPwoOdgDtiFz3qcnGmGZP
77tyFQYb52WdN1qnndUy8rha+YBkPmCwVBQtLenIoQuCvDwKlVj77RNNiYiIZHGh
I30kjPtVNE1MgOnHkJ5WN8VlHFRtvVE+GyFs4XCmBlyXl8d+Fqu4QihHX06xKc0a
r54qkitAoqHbpeZci68ZHhdiOVbcJQoK2XcqzQxvdIhL3Bq11FhdXC9pJf7l5SSG
f0N9ccqZqwXdyW6SBDp/AV0Z4mcBe+2Z8Q0BT+ABFx+xQ7k8ZlJ6SMkOa9NTl2Pp
FzuDWqT2BT8B+tmOdU2Ry3aHVcAa6gZ9I9TC+Z2WdR6gvADuBPUr2YO3r26QCQAy
HPWa5XWiRCthQxHp/2ySurdaEziNcSr2NIachZ1of3Na9eJUKuMTmouAJ7wtKPF0
rbzSg6WaZK4DdfLEPdUf/uTntQTY5N7ROPySsPxBm0XyNGfZGdG9uuzclnju3N2i
BEroiFGVF0Z+2LDaI6C7pgYSZhg6UePmTEeOPv8P7dde7uC1vrgjkQ7moXmlWPV7
7Cm8LUMBjsA3q3CqneQQp8iqVNA/NkexlBZ9MXm/S6mOhvDFPcLSspSok7wI0cng
S1e7KNtEO8ShBWx4L3bS+Sf7iCAj4C16S0oFYNRZUFBG/SzT5j9EVCOGYbTXm57p
GQaCJS5oVbJGlxdYKlqTsmQT/FHddPciDO5oCEm9dyW0ZaoVJ0HtkK9CboQRQw2Y
B/8x4K7hrc/YZ/L69UFKBozXgm2NoqQRRVS8ZG9FTm8BYN3YFPWTxWR6RS974C67
Nz0gOGQ2hn6df2F7dfE9BQhrbmqVZZcbd2ces5pyFlllFEhR1R8TZHwNoy+PGY9U
d5Hrphlozw8MsxYGmxnXgauEn1O/j3pBjoUOY4L7xmSEumLt8w20KA8ZXiDO/pSp
wc9knkwOlrseRAAmCZCFGWmfXmn5zNLRfWDkujcKorzsScdtDueyLLQ5W6BGNp8j
5Nb6IL7C9YYwC1UWkrrlY7u1V2lh1UcOGN6WzkWMhu27xy2bu1Wg06QVwLmI7AcQ
Kw3BnCr0Q+B8Y99x1fnQdd5Glru2LC7E70H3G7pp+YgzsewEVSxyHahvQu3Z0fkg
2pHDmjUE0VDvCSyi8Qj9M8GnA1ozSAWDbm0oW6XIoIXjjYsn1CWseB+SA0b6DWRf
lwvEOk08aAZh3xbzaVdGr4IzKoxATLKuv7VObHzaOfuAnC/feMuSSQDowPbtgnqf
3DTmWDo1nYBQ0s+AjX31lDTcTip2gRbdrR1EARRFe4SshPbrP9xzsRwNapN75s3Q
+TbVApAFmfXUCcV8qpA7AmgCE8qGea7NaGSmTaKLh2UKVp/jo41DhhVkTvy1RfEj
AXUVGuhNCl/SfIrVXlUu/p3xEpYl/TOXySLMKwwphZbHabspsh0bn+VNEBdHvfW6
mtHDxw/ASoJhxwaquR3ep/XX9UiheKtty14PYYGDfWz08tlXQZlsTwikgzyGw8s6
3CzzJsfjr3KDmJiLdY1TDLGYQloF5MDyvWXr+UJfD142UrKRDYVeZGW5NJgEIp/0
DinKwUPaOQkXNbSklcU2p3+VJAel7CDX6Zw43x4HHRyQg3k6YPDkMHp/zp13vV1V
/1Nd9cYYlnlCfhjeN5mE9tKSPFV0D8x85iDASoRb7A5au/8gjnSnBpb1RETjqaSH
ZWletDqXiPSo8m7CLIZFO9PKnM2sCGrNv0hNtB7xkAyZG2JejUbit9NbpTNOaH1f
Hn6bchVBi3Uqjl+0l7VkbaRcvnRkwDk+KHPjmk+XtdJdBqmTNeVm/RB1N1y0J0jL
9kUd1/KFm4IRdp5R3tNzyEt+KwAfXrI3T9qbMZ0p2iNUcYKrKNDgAUC1zh8zEHDP
+b4wj7usMRAQ6JScjFjIlbvykTuLr6idw5yjReRVWXznOT+OZMIYw9ODUMmHwfmg
mQCgQRbNJ5J/N9GutkPayRaitOf09PfyXCnMMbzwGmKW85R7h9uxU5KoN9tfwyCK
RH215NysLi9Ni/WM+RH8E1ZWhCuXHSs3NL+JkKySbJ+dmSB+sIs4TmDYvMJPX417
/INQrZP9XUxPf+jE3npolFHJ/iFKmyfT8QUD8go8QfTr/VMRUUGkbKS9KjOgmRmc
5q/mZYygVbv3CNBNtfmwluVCZ+onfVEZzE3CAa5T74dP7vj6iMS8a5SNpmmpvyX+
7Y0svAIuOv3lbIU3/lcA64rAfWmQyokrE5dlf4xYh6ckVkBNEgSW7xBpaiccGDVj
qMYyLK6pbfifI+MiHKqVfKgRjY/YFOY3dAwIrnfWFNUVek9xMUcYXZLcldpk7B6L
C/ORRM9b/YmC8hDYERHsT8HR9RP7zCiHxmWBCnwCjh9BILTO+R+wn6OgxEpQq3m7
HDm5sYIINo7kvD/3zYl05nxZdj6bPhksd+2F0JSY5DKDGUBA+I/5vBYz/z83ly2N
fPMXWATVekuf51BZ+ljVaFRiNfkZ7VXOaVafQzCBAk8wAcMNDvK5loGAVNZmkDlf
VM+fH6pgMl5xKyEVmb0Uw6cVjXo8ldfjT2ByfhT8K+0TzvnxfhoZeDSOu7sxJ6Z3
+qE5BWF+b/uwd3NerRsU9LJjgqa2ig9sZvKbPO6ZBBY4Mx1H1mxnlF/Tgsj3UWzX
7+RYyLpz+LU3UBUJ7s4S0R9jZQuWc5nPk85KN92MVR0XUrfILKzEuYSgNMLhThLy
K8syqEF6G2VSGhLC29xIjYSPohWsRsjP0SSjQuudcGJP130p8JM8eJr6MGfMtKuJ
h1xwEotwkvdhppnmxq4G+zwuMat8ahjqy6SzKxCcE0NFvOv0bT2CBaCzku3yvBBz
neLwvmfGSWJGV75oq3NiCn2vuo9Ch16wH16fQXu7tWjzYB2EyfXrAaIGV6+0y4fg
yZOah5VN8iHx9ETuM1MmsLTFAdrT9EL4CY7dAKF2HS9vc3eC2lDkDT4dd6qRevs0
jaF48VqJCP5b2pC6KXkcBwxY38EMvuCO7t1pGPE05kpi84vIMEmFwnABMg7i8Xla
EV3uj4CwRzWQTJ7BPt13I8LMaNUi4K6qeVjQq3uQLxnx61EorwZhIxLXVc88LGFP
c2c2J8bFEXbnj31IseGKoLSFzobE4itOUtRryTljEL5lZOFwVoLcAP8v+MMPa3PY
m+3aswk9rljg7Nje2tlQRNXOTU7qqaN1NFOePxQ5C3j8n599e2bQQbZSmgpaxT1X
ucmoo2F2sc9CpTMmwth+GNIJNvUat+HhOf7NodBHuCUfYqFwUIvW481OTCBg03Zk
HBmYoXYubalmm5mFWsddbJpxeZDHogp+LVwFtRd1UY3U4DghYiTDZgcAmVPuQ5fH
mfTP/niK0/7xNsT/jjsSD5UpCEqVZ2HNtU18nBlnhSsGe+jS/VrS1A5Xulssu4f7
pXGoqof1uXGe9xXhBupHCksrCXCaIBPpGEfextTb5kpsrbNaBsJ4lDQ3ZVWQnPF0
ktqr0TFnmr0vjAWo8Nq9W0ZJAoFzpzUGJfxlmkB0kZLfLX+2k1zrQOEBOILWvrdA
Q7npeXuuz3AjR/hYF2l7OCEopIvw6l65ZeqBvt8qpGQSDQXFF+BlkeII/uA+xTzF
QE+mvQ0HM8WjQdJlC9pV+EKnoliBcsYxHPOAxsn4NVtewF7uxgI3x9kEvBN60ljG
J5DCFA86Ik9V/W80WE2rnP9vr8UnKyZePhKGRSyqapcuZcuZ15yMDSVVt5JzWWAw
IOTfMGhahDvnmsVPDT3KIPe2CbNWKgHDJJYcm/+/jtPn1jobxzqw0ThQSfhBGiHD
FvTt+2fNScQ3qC3ozCNFO/0Ui3raFztNnnrQGAjyNzwwQrZggY5ysfwXwBlO6ElN
OP9rujiubA4mUvrfhc0msiA64PU675ojTafjKRswFVZFImdFz6y6YNOwEe8YUFiN
xb4JdZHbZCk3H1p9YXqLl9q+reZvTRCVhMq8byZdnyZOeXV1DteFkJxTGGIvzgb3
rovQ6p2MdrXnN8ikSw7btAIVecm3myxGALv8dbjctl3+rH9Mt3yXsqeXuaHQA9sp
uoBLwhz6/2OC8O0St7IvNHCZieR3F9D8wfxBYQtbjAPH/tKtrVMiykNl88i5Zszu
weETZW33canOh5AP/TVHUS26sMQWrxxn3tx2fKaTPLt6YJSOPsNr9qG9+5RfMkMO
i2b9Dwk8zAB8xLVLzEtjZlsZTLVmGNnlC28aYpzEBkugVsEpsU0TR0HsGx68t9/A
PgGjY1G12ezHJVf3oT//Gwh/dwjB2x1YtKYJzIurbXfZWijsA6R8RlNxKzXLEw/3
VCjZurE+0k8DUAqACuQ9Rm3LxJL4YMiv4dcCvR/J+wRrpnifCAGmw4oTcqV+VCxP
fafOQVfcUKeJP3wiIXdMJVsIQCh6aTvZL3d0DkM6aPX8EiY3NDaUdU3OAkNh+vBY
81Lo8VR3TuSLJW8oHyRZtXqf9So/+eo3gj24RDrW+VkUHh6rMxVnIwG13zPe5KMp
v8+jNDQZZ2xESNYkT1B1XKAjiML4rsIKOo3Qo6E82SfmcA19nF0Kz5gm3AkyRgE8
qgaaRNMZnO8IQAkH0knOraK4e7p4q2mRt+fgubk1HUUGl+xLz4LpvhnhZkov3znB
irTA4AS+J0FrQB+plyk0/7umD2WVwnZlbcPeBLHFZ2ueBAsplhHrhilNOjnI8mJM
Y3SMfhtGITlOfZTS2G/ntj0BNrB9X4BNQM+Ew1/05xV0anLQ+1vfkC7ojPPVKEws
Mt0AmMfVwWHaT1JPCa6CyvvPI69Zp07+u3r/XCYvBHk+PzzrE5hQsYBhdpf6dXVv
TGTbWXGIh9Fg4Uqg+6IY6sSFCvEKJolrMT8TrJbYmcs4UbH8VclSnGXsC6ElDNrY
97RazBDD+ksxtZeSy7prCHj/2hSd0VmxO1dbvXC4XI01OyiZLmpr4JP4ajNWwTCN
FnqCAWcYvv4TncRRw0ED4A9eJm01ERkJjDyJ8ft/veEP12enkBBFLRI+bVo2STGx
VPU0AFFSrTQoewfhrxkFRpmKYgmoU2fk/0SsIVYQqjriCMKbI5YC9kNvRKqSGSE/
m2x6cKI42YXpBo8t7D85M1N9VhCa15bTS6I4e+kfA+mSBclAY+kT5EBxAWyMMu32
4ZpGIDfpKGLmVz/LFv4lmGeZZnPNtNYHUl6FNaKarGod11Cpkt2skSO4UN6lDqpF
XCzU0tu1faotcaVb4EM6fCVhqj7nWzpDFiee1WS0ScXseLcd08ibL78NfvBr3Tye
anCgTpcbjScmQOj35MxMykxG6ul0ywzkGWcKNa6PrDCqhRuszHgIHwM9N967EupU
Z8hyIb3oq7xRtF8u1SL3KQgFCP/3kteL/oj+aJqugEGV93U9KTiUQhJmPGCFLJj4
pu7YtfYFRsWhOD/PitL0W+9VHBZR7El/wdRNbamMXUG1/hdgjQe2o9cJdZBAeJdC
Gal5j+bZD5qnZ2kYGQJQN7s8BMloaG1Xm24K8kNxG5FtmFreApxXu/53iHIvZ8Jf
u7Z/0p7VW3ALbN/+eFLNEbHt0PcrzrzzzG9slk+pbXMIBdaWmbOJa/Hup0yaconh
YYoFTYjU5XaurWXuOmJc0m50m8FbPwW5Y0YHp7cb6mvbdeQoxAq8lFZ6TGVn6CIP
jR+cSRpQdFXFWa9z/y87d159uVyxztFgY6ObeFNdHV1d4DtnPI0BJeuWM+V/eA3/
vEg6878cVYYkGKMttpYkAlZp7sx/x8vtTLpWaw1qfGS1fKggFpcX0mJgc0y3RxB1
HjDomYlAfAHBWaqRCMnG/Gy2zhOzt1ySsOFi8BbYX1P5955B2v10fvoNvlZxM3ds
reofxhbst/k6hoR0JKoL5Lp2/wgEHRPb1gPupALWBvreuqazUEzo7rbu8/Y7PnEt
eXQjGsSNopUpUZhqBBqUsZdaxsk2zzY3qPukvyU58Y8yey0ayOuGHdLN6ZBOZScV
2oysjC1Rsod7trKotWshUVdY3owjUycpzoZgE5LZkKZtRSkwpCS7g1AohmgHMGsW
ATzZhau2NNvAIMqKrFZ4BGHBKXSkagcKfwvL5cVV0rD63yMl2sQF6StGW8fytww1
KylCMAozW8ovvTjGgq/ihZNuJvxfUVVWrBpvP/+yPqXljxPrFcC5GaXoXe3BSbCp
wsN+vil1FeFg8BfYvIzdUBfXbt2FAw+/OAR4iK0Alm7JOJ1uUWy19ZaIoqlgtmYj
3LevZp2gWABNvNRw27Cz0ekT/+9iBuk86kd52L0nlNsr++3nIAr7Qysx1f0dCm+3
/jztQIi5eS0fWOZbBgZseKkElaXOSNPWhyaJx6eFkYLH4URnCGXc5Tg8uwDca9bE
aJAC5K3Afxm1o2DBUw+y4awMOpWe8ZSZkj/wL3kIBIm1IC+7jXUZomHyZmJvxpKV
OWS8+Gl13899g2emvfJO58GQiMX8ZExw79or8cDvE5dZsXXvRy8pCemm1UJkyppr
cF4yCBG28Yb63NioYYhZXLM7ieAr6yU9SH/fgv2TgxWbG2pgpJtrJoPMqsU/wsoX
93caxMIUU0Sjqlg4Q9ifTw0m3LTJ5b6cVLToPolBRHF1tX4B1gdDkfOA29uYjpv9
dfSxsMlboV/9vcsozZJRtGSpUp3Cz0jV3NoDutYFNtSY+MOc8QPAAIXTSRRe2YQN
BUYhMUBgH8Q80e6wHD08ylErUviVL5rOtPHT/hxP6YsJJwnRWApYx6QNwrN3f3UR
UE5uDVLFq6QqtfREbDDwl1LFOLZ/ZfePdydtdFO3E8uO0o7emGLY9dLUl0rkZ1Li
bF6MUYC+MGuNFxKPXT61aCG4FRLIkyUt6PtxqWFGzKQ4Su/5PvRzEkYvuMNDzYzp
KTZpTtmfQPtPgQ3aqOlO0JR55ksdgFYN2wR19NpvQrWK/DbgKL/pashYd7+QWArw
cMtbL61WWkLSyjZLn2dGsVZ4eIpzW6hl5dnA7oAYMP80Wqk+ZPuS5yqOXWYu3i3V
Kk80w0vHO0JXDuYmrYrefQW58ih9f8XFIq2jsx6pM2E5qu5qV1Vx4+2mOuDsTgc7
APZwulghcWyLyfYCc71AZa4ZVnCOzkJoj2py5LWCbl92iFGuEzTNfFxoFh0KDQ4+
HkZuQiZiw8V1GJwdLraGgHE9c0OvhKKj8mJBFKtjyZcQEnKDlJfurj1fsTU92D0Z
xLnIAq1EeswQ4I/gWEw68peJKZIusnPy78Ork/9AIUYAXFGqiiNPJBSuCpicOByM
XFb0r1Sf1bTpytKaVcJFrRK70KRMXE9QYKVroEZInioB5RvQ0tgRH8PnDs1j/pm2
mpZ+nD8tjez60PSxSDbAFX9dq0rGeOD9dejIm9o6NpbZ6QD60OZmDxgidM8yGU6o
6/7dOrd/Nq75T7s6cI5nsEt1NXjJ2zAsREdLoKobd11Rrs39O1vMK3ZHv+hapFZx
GV73h/lOX8tz25PGvQCQJu/8eQgpVmHTYHuQHYMlDNNY4ZIAzv90EjxndO+tEvnJ
Meoga3zzB1poixGFcnwY/kEsx6yQMmjNdHF/ds3rLEWUV7wHbpMpIyzUdDJVXdUZ
yEz+3gp45moc9op8ch/4nEzPQ0wJfJ6oAwg/+SGmDIOED7N/9brQN3F3BcE5TBQ9
JgS/vFL/tRZ/utpBL+MWfE1AqHdAGhjQ6xHDZfzT1Pn1IstUffOqrQNeUs/lmcsB
avasI3ZpAhbOjRq/L1F5BXKLzZiUT5DJ7ANMHwGmsyY3suEtLby/sRGKvQt7SHWu
u7iZljukaJflSiSa5QwoYblrhfx+JsUr/C1OdfD1x/fDy/ZL9+vAcQd+h4a5rDoT
7NbxJBDbvVTVN25zGtaLDrFV/kUIb0m7Mll7bWFs+HAtihJR4r5hDZ9prToqInc8
yy2VX5gyc4E+km5Jv4YXFJivgYys36gYP/YrORL6FnufUiC1d8JcTxfa3jTjivJQ
vJz9ZN0cEMwry+W3SaM3k2kjJgUnj3tCKaxoCrMGbWuXYICzATXv7Eyih20QpfGg
tc3jWzYWfIaoItqo6k8TyrlalKAcDtEG64LfANB7jMcs+ZZmc1O5cBnzc+7/fxoT
9gK4FLnOfAQAVCoMhzbdcHaO9WhSx0D7JcMKXEP8KP5/HIyAGoIMNQ75NV+i0OUR
2bv74OBTG4R7Rl1s/2ern/osoRwmyEwDnL7BbMWZa32QADAP4utrnejRqpVGTXwz
p9wCinSvbs16lPBUfA5vLCZ1xRBa6pp3NZdpTdCBERcDWTgUIzT3J0+dqAtPmlXF
kg9Vc7GZAx3K/6vB0FaZMGovakRrSKmjQV6Y7/+HwIU8Dto3gJ0xPL0Ww1v2Yw4g
+ovO5B6EnhbLAE6q0LLBXFOooExSauA4Hnmm4dZugtoKTCjBQ8tXomewFJ+rwDty
sqWgYVjD2uO0RjbbnCS/tTh2N5GBwS35tWmZVnq7j7crK1nf6bptT6/aXOoRRhuO
0A+L0D195iCFtP0oMIREIKDcgTez/x3SOC8nCDg0szFfgFsM+SKddUJXF+hHkQRL
/Cz/7Zzwkuoe83TyGjC/lOqla3Re1eMdG+hGPDwMLRgFZxHsTwZK7M6i7jatLRkM
JAj8nEgj7Rz9oCdiJcjvZmGHh7VMn016+TUB7WUhHxcfRDKVoIIgMuz4I7Nte1OU
7v2ANMpHPlZAu0qMpvMzS7m1k0P6UDYxNid8dWAxLQNU1eOGAVONPngA8qAMMFSk
V+AsV7F9nqZRlfwFqL/XtZyxPjiX8RuDccLvocPYozcetd1Utx6XjHhLJRsECmF/
SWKmDg527PTOwdvRGIeo9cGB+ty/JUJ9aloZqDjWQ6lwvzRFMl8sqZ3eJorNZZc4
YYHkDCGx1eyGNBvxw/Am4+SM8sCNLuUxPOINJDn5RFEvg6zut9ZPd/dD/9z53vyB
gmtH3IxgpLB14qcHWRT+kZIHxTeiRXeq7+QksZUoulK/ATwJjTZcse6LB6GPQSsI
KZBrpoDgsErrVkxHuB/mHzAnUyttnSy0LazZWRZYsO5M/2D4I0E2yPpXgww+lYj3
w3qN+kxPX0/D87dbyruT2kkcnMwj5R7sI2cEZkQQOQAwXg61/is9KMfQxRCnCehV
X8APVseo7o8McBw+BckaooB30Dknx06QqIQ2HlgN4hMOxossb7Ir//37rQaAyPwU
+0g1zJhBgpD58vwJQAuzfm3pdMgp4DJeu3PNEFHasFQELiD7bcXInTFALiiR7PGX
l2LkOs4oCDsMg0wn1jcdFzL0u/tXuLVCYGuhxE1/phsDFFiHxyKtL/OJgM/Bv+jR
MK2EcEKSlb4r+TVNnG1AaGoizM4xZ55lN+eaT92haVFMyHwJQyz3YeP2fl11iMSD
nedusQWozQ2/wTRSnGBpr4U6K8FIQtvCmTXCvpOjvvVncPEC8DSnviOWnEXwCogX
iaQ1Z8tiiJ0vdQXBCacgOFVW4xNG7c5vUN8/mmSI8ySPGHq4VlvAvWvqmJDsPBGN
csjRHrykCeNbkAkmhtG8UHWpMIRlSeENennpU5MIiom5I8dJLctb0T2WCRs7xJE9
2NGFK9IkGzo0sm1TziMJAGepLkw+FT6EmNRASH/LmiuZKATljBrmdmbg4jzCPKzF
RaguGJcmYaXsyByCMDAwcOtngWBh9M8+F/tPHoge5fClhoKQon7goMVGi+mTRZCm
Q+bGLkI6gMh/eMznDFLYDfBOyc/Q1UWlUrvmMsqH/NFe21+9pwEUqkGiQaNJfvxF
i/9PV+6V2E8Eqtu7zGJejm6PT1DDSsL6txIh2HmW9WbJ2CbyfNP5ckcWc7sW1qqK
VyR+UjDxaENdk9HI+nsacJo1hwJovD/WfA1V3iOARXfKdjIrZfjvijZTO5pqomi7
O7xQPAGZ3Elt2m/+ctHAUNRNIGO1Hwm30MIz6RboVYDPGYDlhKfnrXPd4atitusB
Pu82RGmNratRw0WjHaYFASwyQDvCjch8jvyewmQDTTAyZc3s9AjRP/VEVyspprzX
tp5qJp3k6TXtjw3zJLUeDivy1OjyRZs0B9+yzE9uhHp4WarxKvHqghNYl1RhCW9F
ctsrB3bFJM7iqHW0iS6rmb8h7CvLA5kr+8C2ALvwO+hvbD+bQuTssj01ow1sJ27u
uyaPBDWX9CXQRCQwJJyx2Pxfmvic4ammYARHsB0AOLrXXtBa25gxM2GkoX9OEFxt
cY5asZVNIlQEWqvd//qfTcrj2EOdq3UNUV9S+9q628Kmk7xbCFSPnYocd/OsOmD0
l7IGLgCPNtB8f3aGXW/xRvslLL/fCAdisLx3sI+o/5Z7wssyZE4KwSGeQ8Ed2yyE
64JTJ5YXsyekCheXMAPKVZ2DB1t5pCP5Rm/3H3e520V+AORG1q76zyWRrNnZk/V6
RzlDxIIqpzEmIecTh5TD7ci1QHqjdOZniPd6tgFs94V/HVKI+BwV/xgoaBiD67PX
sWHa67HWLWOASkaNtrrKPaheB4LxXmK84jwbkadNFeVsbAchS3HlMUyXGDmPIM6z
ZHDVJK/OI8+zitqC6hfG7tJW8oWywOrw1vsG1h9RakHhkr6uQx266tAIygVKh0h7
IteXKxfCPzm2Y6kU05JystpulngwIWLY/0WxzoXZUsj6iajcHiEHR72qmgP40MfQ
cHEpOngp0AHWkCq551exfnDgPIoMnq7LxsWChZ79jO3CYG3S8f1AltzI7923bjrO
GeW78MhO4wx+P+BzOGxA+1XBqT6ZsqFPc3D6jWfCi7X2gUVeiLAbYfomEYBPA5F5
SDULLUZ5f8Da3ZKaTLD02wzlZtHsNkn1D5oqC2kh9BZ4hO/zzmZsnTvYgexd/I1U
i02ggHj4JHlV4DzvC26wHS9bWQOWpuLq30uLk+gttvKl4DGYGwXwLHlxpbkt8Wli
NDupBYYWri7XoZ+4IpBdgqLvP8yRW9o0VXMGmpcSoySwaUR474v0yHLQIYTaO4a5
a2LL/q7n4BNd4S294niwFz+NDZ7y9fVpnAd3rTiA8GtfLfE+cS9dcQ9u+X/ZR4qG
inkEnPD+YB6hjMOu+J/tK4IGrzWkKNm6cT623uMXH2eaaV220mmdoY6papKbTvAG
4KYjvKJ5EtVT9XvShvleZyuLQOXdDRPxiOdrJHTV85LNL518oALvxP/TCP4Gygbh
2esyFtk1aJHBXFzIoWeg3CVaypiRkZFKC9upcLrULQD70Y+Z+pDPsJdeIWh9D5Hn
uY2LMDtePbo5XgWPKD++2FwkAqW00Gpi5f6ouGojogMhsu9BPCpCGhUNGzoCDpOm
9sv5IIfNjRv65hphNykDrWGgsNA4BhsP5mwPZuvBPoBPCU9ad6W9ZTJjwn4lhO9B
bv0J9pDbdPR/DZd/d7gqsTe6ptkfkTLoWyaP53Z0Ag25GmHeF0zf/vfJLUQZjD0b
IW99xsfEu207O2vxAMpFoC1S93rreVvtDcs5uFN2amW/MgihnYonj68kBGo7L+4d
Sud9TADu3C/tZW4WA0cLQYTFxNUlZo7Oht1HAo6YbdVeCRDse8d78NqBrrGr5b9P
JN2IELoRk21PRcm9AtIcEMAIB0qTcOz03X9z6MO6yCuBzm3gpaKpe8/as+q6VkPF
Xrj5uMlGtfoixhuwCXbvzNS0pkUXiVNbQGji5P+HRdFAFo8oQB7yjlnPPEVJ5ixX
eAsxVpuyeqqCNbpitB1BL/GCv7r10evQ6EmPaaikDy8QN+0AVNFOlLaNqTBnhcQw
8UIcuorXiemaXv781vELfW7lUfXxcaVxi4B2MyMuxUH3MWwFTQIjiNcZfHSxy05q
wRI/LVDTgQbfxGuOznuq6sqAP8EJz5xYlnTKpKJTjvmtj3ccxRqRCYjCfU83n1ZN
+jcxlcw7AaTbBYeqZ22jqsT7APT2AUcrP+RTEcl7bgACHoJ1CFXKtHaP/COPHZgy
nryhQMkmzP4XvuGjKcLlVHuh9ws34DcakRIfCx1DotjQnPNXF3fVnrheQ4kJA9up
NWyS8U1OpueUfE5lxcy9jywwEWYTrl4SUQoyxF1yVJU74RKsnrIyr11yjhgPilWw
+tJxPxpFkRWmZ1G4z6GEdv+UvXcEDh+3NaQbV+iQ6vTVuMUD/LPbgvc/p091uGT6
4SRkZWSiuWugnmrXKNQHFHB43G3ORMgGh+4y0sUfUZlr+/VB46trbPnCzaGyW/f5
B+a1+OL2h9IfTEQrbQf0RNjc9Jjqd+dlMY1xbraYKKtm9q+U1DhWITfB9PZYbdPN
aUkI9ZCa2nXHnPw9RLKNoTR8uRGeR9dQkPP7DSfb2HHM5k9aWStHag7TBleME992
nfmkqSt1kIj21Q8EqtVUr1BJqqw4yjA5fQsJVppLc3G9LTjPPbBVn0CJMb17wsEk
DXdgdBlR/o4iNiuvSB8dqEGC0pXbRfwFuaP8z1PL+/J+wd2wgpoOkvgN0eN0apBr
41q49wtRBDMovHTwkeisWbg5YhUgHEDmwZ1/nBD8aXb677QVV1AcoJQyHUVSGMm8
XefEXMu1Pwf9/XxeLLzWn9+bmtnL9If3MID6XtbP0cwtfNmSQ7tGHGe7hL1sdLfe
uT5vfeG+7RNS3pe6Qpn/eV/RzPXRAK8O0j5XRzdVAt/FntZtdH3Hs9BQGi51dvhW
cexXAAuokez34P6W6wStOOBAaHObi1Mf5DWt6PBa9AWw3RBk5lme3fK+E7ivZocm
l7yvSESYE+NKgZMcD2QTGu/MqOCa5WAoLFRUaKniM+uF1sTURBU29Cg8+0LWSEcr
lrwr1AepXpgDQFIsFGCszWtUT5ZMZ/PeMsRhb0uuc+8QiQ+0Q7/G8fZrt8Dscr0j
Qwbul0Duw/w8mWcyBUFjpReuJDyLmAgZXIMlX7wLhouk9fO9n82oKPN82gXVUbuA
8N5QHYiRxxloqa64vEEq/saQVAVHtlaWBi7Poe/zyBoOHh9y+76bxNAJPujJV1Ps
zdvgEk1yx81hfZUrWbMuUOSmCbrjb98eKNCWBMykyXA3sgjFUoW4uZtVQeJeKXBH
qTapVuThG+/SSw5b2cZxHy1wSQmIRVDWi+/sRHSk0GP47I/rKbI7zKPjP23JEypW
UeImE4CnC3sQ+d72mvnLACNN36uKj1aZe9Wh/m88wRx32whgB23VUWeQ2q5p8RPn
mA0V8vjPcPxbB/mGgodPv6oZ7OIU5DCJTzV+ll8Sd64Ud85c8UBQsV1JxVrmYbe2
M4J6owxK1lRpIZUBaT4f6pP7q6j/IYrv3OK6ZmPB6VdFAOSk9hpm3FigaLypeNgg
NkV44c5BS6r6EccC/vioH3AURfaxEQ7N6sVK571hoszGaC1FCk/vUP+dnclWuXEs
WUsho3IMd5wp9mbd6AICaOqoCsw2c19Qrd2LO4LjCYDhiDAeV7RgYNccgfZgR1v0
O0/CKSbpBFfm8BfIBfnCa+By7VSZXbqIAT5Ym4XLxkOyX4cf9krD6F7eNpwd5sXl
0S4WoTmfMfXEbXl/OyQ/suscsEsN5w/qbHok6lwOd9Erqc4uITqstUGsaKrXGJ7c
8uVt1699MT/kc+HIMI0kHduCtqgHwZ41UQlxlMe4//c7qpKq5oAUPpwZW2bZTxVq
uM/jJqpjy4pE/tJS023+jM0f+ARWg2Ls2YGaNK9Wb8WI80meh6CfRqARe4OBfM2n
O9scnbvIDVxRZSzNKnZSNqNY3C22fPH+Ndn6ShRm1WJt20HkdPFnqf2hgb419m0T
Ei34Z2oWxyz2lDxe8d6vL7VPd0zh3Dnw+qTfZy8iQfe5OcZA+XmtGFVpiUnYfJoH
4Amt3sJPBz6Ffx+9CioeO6APndQQ3S/SUA0kh73mXxeQDhqjDELiliyu6OOksl/2
aPp2Wpw8iEyXEuFTHxTUqUKkKihTpGRuu/TAd8TVwXBNgRVFApWiBmxg9aqcZWNP
/pd8/xjz1YU5siExQ73xUrwHRY93cH6nCw8lFmxP+6OA7zHmqzlgEnF1Puy4Hh1U
grK3Ox9mPfIDDifs7muZAYxYQx8nA8Ca2umIyU+ai0zGZxjRIsTwyNao8MpYeNQ8
wDJxsb1lFZ0rj/OB/baIzulOMRF9kTaivoNt6V4GFAWwT3SJ1UnYscyARxXUkaJ+
yNzEoZNiB5+5ODssJy9LOCQgJDAaAeSwW9+iONrLCUi4wJZIAq5Gaz0sSICSG28x
I3WfmbANUyQG082dtrZ08qsAj/qsPMYzI/6uHhxUPkQUr7TFBPfoK6wkPq6axyDd
C2KD3mW5AjDaWNUTRH9r780eHkxYIlaa5xQJMYnK2v0Dzgp1wdmp/J6OLlhq9M3j
nKDnBbZFqtn40mBfjpetkbVVK56Okee6lXpYG+HkiKhH+H5+LE6WwrKJPpSayyvf
+dzge8qfqhKE+JSYJ7vlfjuyE8VnQDwt5vHXdUBDNMBC4PB/ZcgpzdZetIVCvDFR
A2MEHs5NR/XEHQaAQ56BPTz6Nx+SGUnycrJLFsBvadxiSFN7tlJEyaASoW1ocfj1
vFtA8A0YwMO2nBJKXUdCtqvCHimTD1F5iWzBP/pnOWpnYc0fcSWThveXBs7iGUAK
JH5NfnczbK8YZ4PzejvsIWft+YhBv6KwLOiOqbALJsvAc32thawPmbtHD15Oy6vF
byRV1nPzkYefRpKGuYWY6cVH/ULu4yKvlxY5VUjZ4jLbjFSv9Qq/tEMRQXyZLRp4
ISFR7kXANew1JwYN0NupMmT6Ozashk9PU9fFlSnD1qiIlQUQ+Rr5TxralbDY764v
sapIO9YBaR02o4VzgrRP6Qf8HTueQqKY4Srd4/Hy3Y1387YMCCd6gXcvFImke8g9
pUKa2G4dJDzSA/NDi99H+wO23alpk5Xu2VbNqKO7z3HqMjyoEEK1knrpspauUk9x
Ek4hOoIWl+k61IhNnVgnl5pL3kCAuJPoFlEr2wr3Fo/jJ9xOM6MhnZmRvTYRc824
ObH8VLIQlV5/zwYwOstdsGbNpUrzkdzH2+eADyFsCIfP8TvDsbzEYcLEDted1NCU
p2LoeW5r3pkHf8JMoanzzZ1VEnVsinKMGPk3rhFdHJgYIQRHekCRw5bToWiezVV0
Or7+vXK3mXSoApyREUOF3N/jDiLBc6WA4rN0gB5bghF1TF6MeuHKB6B0nfKIgWS4
am8Be4/UkefQNar3obo5HwjWeVBlhTXJ1rAZGG2EAopUlFOdaDsKWvrmGBOzun7+
dlS5ygcgfVSutKgVgvkuenWEtcVaQbgcwNARh5xe4pW9mwLJyvjod9g+dSvvg7dg
XG7XzskB4CPVtw/c2sO5EVqQbQhkdQw2vOYCtAR6VOvcIE5lDZ+++F1+PldyidET
zCArdA/euzmwzWcQgiammx4Ayudf/GerjmPBHFi8tpaNXSjCyWNo4HT4pBf4ByCg
+PR3vYXQlod4aC0zfUiwxN6UCFc9i6lvlNhlm8wnloXpHw9Ms+fmCATSqUqOWGhR
CrpxCgB+Nc2CUTT4nrPaYffQELI19F+nLpZ4hqUrgIoixFCu7XKoBbOrBrZJNcXb
8pRR3PclT5ot+bfhfIySV4zkoc4WRWIZeqAeynqNrLbUq+PIzrsPu4X4pzYTiYSY
Sm0Ea4Sz2cVEWDm1qclarP8PSEh0MAXmu1X20BLFPycxK79JPKAbVuhkh2q2X8ns
E07quoCXsTA1r7V3ZvshZC+YPnHRuWnbUk/9Covk2PEQ6Un6npImAg4246bMjPlk
UgPhZ/RZGUEXvWGK5AwlAadB9tIYsU40j6Aph1M8KtpgZM75GpTmC71kWOtAYkcn
fLfSh0KQmf62hJcLCqIxeuOjEVV6+0AfVB79h3WRYn2NvsCcas5iuYkHwistISb0
0faWn3fztFM9ZGvXphuY4a+SMS92AS2XpH2x7rq/Fg/GLshlRYK8rsrCoAhZ3y6x
MpX7zG+7een71NtcyGwhRA+GiN36EWPPgtqoclpOly1a96ilgOzqG9VnRfNbOR1A
cPWSjW8EgXqkKj9ZrwH3Rg105YCESj3g8otCA8z7I3RW8i3iYzzAk8Vs+lW/cPuw
fZp52qrCFQvo2VC+ZmAqtj8FEmQ7uKnKCrz/fw6kvbs7SuKHbcfKHFS+TM7Woo+t
qSLkKIW/YKZw8XGHTwotVS3mqXmZjmKJX2WVxQ6T3JgQLYZ1FnzG0jXf29nu3TIo
R/z3jMw42FKbiccNJcbsOFeE2rTZBsxDGTEQzbdV6UpwFDD6NjwHmiekYxhxQL0u
zeze+iny83cPW2n/DAXlgADNes23FX3j6u4ak8wuv4jiPHXYRw0+W/sjVdbJKjUt
RupjUQ4rnWbdTe94JQkpWvV6Kj/xAiJEU8yhsYoHn+Q2P2ZUTJAleEDj8aOci5+H
Sqd3CQg+AP0m3+SnJyCTSh3rKCPntuFCsYCgzzuI5XjGmKnc7EPPynsMXwHynicV
rJz2zG9OlMK4hxkEXlY1+KqtCAnqBN1lgMJfUWj7tMazzjZAPJLaUe0pZCpEKPF7
xFDk8mlXwH5UR7GWTlmWt1vk/IPcMIiWB7aOLIDUjbOCPDrtGPrSR4NTh0fw30TM
dtCLqF6RldiAlKrgVfFP2odc0hMJk1TsL/A4a2nK8TCa4vt6/E4+052KAQoZOvtu
ZFBm7If/9PxNB6sJBZp+ERuDxxxg3u4cou4jpQkR4T7LJtqtl72MkssIeHnEP/3Y
msDwdTV2R+MoCsypn8gcy6Xl7qSDeSYvZgwRPwLG0nvOM7sYQVn49l/Xe4Ph04dx
XM3K3UzWYbX3pSUuNEMTj6c2dUoilgyQWPDDoxTSOfs9385rsPVvVitE37qpcCtg
XfMRwJ09/E5+0r7Up9t8eVlr80G2dVQZXdl/UiGbLBw4+cMkzts00VsUZAuJ65ES
8J96E03xdy/eR47FZTsEwLDCt4nJg9h0wgiEDvZn8JKpRnR5sOQrDt41btc3JoFd
mHMU8xeNBONC1WgqNktxN3qkkZ4LUriMQOXQY2RDrGCreaV9F0KSTOKerKwAUSyV
vX9Wr6okMxWqeMZvQQO186yyWTqrKJkyeStRi65AHfQeCP2izbl/9hV2fnKgUDOz
mSL5MQEbv9BoROXCBbbPCXiFdYc8yShQlSvJcGq+HpOCkuI6AuCC4SZRKSCIyI7z
aZJksMlWpBxhwVDaqKwmAF3KEuL1pzfaHmXRI4UR5XOLOGqbW0gvMYLaaSWvalti
tZEMqURnoNqZX31AmB5eJItOeXPOrCulvRLXuWV1+qBbeWQjr3Y8UP0x/x5CL5Me
wfPVVuIT7Q33neSCwicqAJz1ojqUlawoWVVA3xoVW0hUIB5ZBrzht8D44smgHL71
wmu+VjCJGySAJquaWdmFTop7TMzcHjapmwvUyRVwTN0HqZPNBdxoP1YyGVDyABAH
sHOYtuh/dDRSjVd2cggmEB9NGDamr2JwDO8tHPOjK1tAfADxnKyNEb/HsN0L9Qud
c+wLWSQkGB3YhPNr5nM0BHl+99eCAxSMIeuHoUYWERwUjNDU+KxmSi7iCFCpStVe
48FC62qDdumusaxR8NpuOFgHT3gcusLIJ3AK1HD9kkWHumNw/gJWTkOYfpnwx0DW
4mnotOTLkvyeJB6lHn4tvdaSwwV20TBNBdCIstUYOEcK93e5aQ2+gzpOoOlyKcvb
8xlgwoe350CQbKufFuIGw76Jxj6+0n+lHAJR+RhDO+oa31m3EMzjs/EfPQ1klwhE
ueTFm+gXB1eAVxaz/3sVkVF9ch5n+fgIa+Uqf8Z1biLn0P7PvK/114CKaG90EXEd
rYOXm7gjAFLEiRVtgyGXiruxnTsKx60h2HIar8E/tFxKfJV4x6qAkKf3cJjb1+Yz
iBgOwA6zquDP8fr3hoBM8/7/2o7+q8YU7kLi6FZVLjNak6CO1PYkIWU375ETh8ze
DK9S0eZyJEjLZNjAtH7amHJZP4i2fUavEjodWJnSLdsb2cRXW09UMu5s3F8YyZmL
5KubB35QHQyU+umBTXLK0Szt7oSG2dc9m3p/B6PMtqnKrIy5D1tl3Iny+qzlSl39
z+VTacsTq5V2qux0g5obx/DXrgfC7zF50v0rM3zbuY4agKh6k7UF5QciPDCTmJZc
evxX+yBjN7ilA3pHZ5j55LDJxHWrIws/L2nEv+KiRT2UOld37lpPQ9FszADa2tk9
kEGuB2cn9TeuxVq4htGAHMmB7agv4jbRz/8MSmDmT/ZcHYNuQbkoZZ0OaSmkJtio
1pKyoGDy95RDUlN6l1Hpd/PRYbK0PNr+h8Qq0WUDpGgm/6DtO4yH0soQW+PMjDFp
ykhKVg09vm+6UlIAfKD3o/zdWyV1gpY2D/BjIGTfxAd3BbSZv07gOblC9Couj+gf
/2Syj75KlThKMDz/+kGomt05pYAa7PSnwUuQYgUM0nADrp62TgAZL9ElalqVfk/h
TClZQE8d/jg6e8zmv9AfnKR/oCdYAbg6CkDHxNETcg36m/0JQbsLSxwjQn/KZXkO
xNTK2aTsmiK+jXqV6SJShvE6GU1pWIVAzO27cHZXoFp0CvBjH85g7YIV8/TMv46U
0H47AMhHaMT3q0FCVUxX0MDpjVaRF/NJYI2aZOdvd/uX6/s0dzPtL16p2b2lTPLN
+ity7Kt1DFm0GH3rjQZT14qiF0SjzcOearXmNcwYldHzhQ/j6TDAUuEJZFsQWYQn
WpIUFF069tKKJk831W5GM4Q16SU5GIvSbk380TsGyxYb4G5IgszJ00MzcY83nYl/
zmKUpUfSCN0iFjf+L9vDJZHqzLnNe0sX9cfI1Ag2tfBuqTrLx/tfkmdore0SPPzL
0zf3dZ9XyLAFhb1jzUhFofZQY4IgGvmus7QHJOcTd7v+3ApW7+nCCGUR1DjXtF9C
F1Xabrg1OxzWjzPxAUz67ai11MIOkykBLpfsG3oA5SLC3nYcDupOOPqbiFTTH2c0
1bcLGhYBSFXmCf82Igojwa/j7EQkINLhlMjGbFLa8ayE2GAltpMExRtj98SQ4/zG
fXI0Yu8DZBhJKF2yBOEHx00I/d8KN5d53BuQrWBErnxIuFaWGh+nYzoVn7fX/f6D
0TpjLj1D3LK703aZCZ6bjZCgUbNJ3JlcxUPysmFNzQH6uUOdnwGEfV9AvuvGJOH/
e8p0mPMk1njivFDYDNcB26nWpbraSY6YK4sy9AzDbz/hl3hjEa5GxSXzqbT9kw1s
zC+3c3CebvoA5h/p29UCHh83bbcZlKFjeti5rbZDGV+AnaLL1PTWpk2SZ6ZlLSVO
x+F0xwAOoh1BkFlpUsZ6CxXOCTzAt109g+OKXBV17es2v3j1YQJmU5wGmgWdYVKK
B2k7KaJoFjx3/wSfeJbt6LVvdCfpwf0d1aQHKTQfEEPnrtSyC6z/VrSQljCFhd+W
pQt+kIRkKlB3pp9hg092RM2eWY38TEZIKh78z1AzSxVYM2ju+w5ggjUPw3dLZnaC
YOZVuaWqEM6fA3Rv6gr7SCw/X1iaNenmk84fX70toBHWtU5gogUN/jwM7yMqDPfN
eGFC4LULNINcSrl3JcuYSSQBq558hkh/tPROGyUtyaPbbBnvQ/UUC6HX0WlRWSFh
cAJD1xuDKTXhl6rikWYwoEHmtmhqtbnfqLAAdJg0/XzzHDDUvE4+bwUgq+ixZatZ
QgdlaMyI0I+5cSwK+NH0e4QcXji9toTptmh0nVo2jczY99+6i8bZugtusotPjebT
398/e1bVetfqCaD/TYFGKtnFww5M3DQ6I5rJeAwyUY0+bKHcRdkuw9/BUEHA2CGE
4gBGbT0u02E15FTBNbgo6PbbmYd6sGWHx7Vf8bKg+HIUELtbsKCf9cL0ohyYKOih
imKJICG79YZZsBA2uCwqWlOt3N7Mp7ezEggnZxhcebuhguO2c1C8blWvW0mTEkBY
gE7g4CcGuzXmQmabxCocGcT+EfYwybzocht+pGOkkVhms/XTkMporE8BVA3m1snd
tABgap46DLMKYis6mVSXERww/UzJm9nitDY76z/EZmwAdEQqNBL1tvTPbcDSFFwA
sKWxOGLXNls89HC2KK861djZmOyyneKZCmJSUAxDcKavwB9KbfclUzWiL2uKPUQc
ml2kWZM5EU2ACi1prMlKpFNBfC4te5fC1etuEOWXD3qnoq7t05Igr0nuP7EtYuAT
3vpwR7wv2sVDaw+qNWW3yHKmPsu+qlR/PS9f0RvNesx4C2JcE1HwhfrwiMCRLsta
L92e9Iit5ixtcM4dw9999gJcRwenIlONrftSz6Jod8qBohXJWoUMAIryQTSgbyQ+
HUMiJ25QFtlz98Kslhyp7FJeeOqZ1g5UlM/JVx0GGleHcmHeRepW1+QbiuV+TnXQ
NRDC2OFwoMtBSY8Sqfa4cjubYPuoYzElAADIIoNKB/9SQBJnvgAWpZBeAe1COC+H
k7M0PK/BhxyiRiXvnpt/ldDDFyBYMebXgt1D0AzBxrUWJaBjbX/M68yzKr1XsF9L
Pa60y/5+TIZHwEOiA74bMq0mMgVvxrdmoZTG5Sj9nTKQfuz6kteLN6PbwHGrzCwC
v0nG45HIUrB7Y1K/Tu4CSa2QMcNCfKhqJPfNcfnm7B1QZplMpoyRpSSikc9MPBiI
w6qT5nYAns9aCgAp71ywqTWVQKcmwsMzX/BdpBp/7dGiQhxwgaj5HkHSSvQWGQ/w
MfGJoVA0rliOA7uoNiCsJqxxK4C7mscXfJewp2aazPxyj1r6qQg0AjrbYPoTUtSv
CPSUkPl/hOIrjWcgALjraBYFLHyxlfp9nSvKM+sC+KW0lpGzxSE+PXWFM9hBMx2K
ZoelzIue8pAeEactdDHtQpZlNI7SHtXsKnDzMR59mh88KFILP02dYa2ZHsFOcaNh
+31YZMyA6Y8coFL5Qi49GYwUhWqh5pZnKpTzkhK9Sm0o+dXGx1q0QOpBB4jUUOQL
wFY7AtJISMMsIAcsjuHWbRkTPo4u/rR7LGcQ9HkINzAeJnG3KTvdon48R5uhlPyG
fLX2qwcwnHcLguorlIT2SchwWHjxN7KhucDIl/8jMBWlOM+JT5LnNJckkuknG3D5
Q4YVlvNuxuz9EOsu1oIw6cU/mUHmdWRq7ivJ4WHiZEGSVd6l9wTINhiffqZvIcBE
2jFUxagaqG6a4gHSf3yvpX4nkzW0GSuNT9t9fLxpgsO2+1MNhUm1l/VgxtSoPcAN
X9hcagHXs7l9gBUiaTEm5q84JIp7wEI0V6KKq16jXZi0LQKHWLOcydHyORBd4OoP
RNaqBYdttw5dNu0pMJKjznz9MJJsSrElaE71HX2fRPaccUoeq3hsDw2YFmobFjzl
3XnsVENM96YAMMmxbnue8uvop8QL+jzgblnDWK0xgMdUQDir+lSppWok6jQyJbIw
g1bUSf41hw8kvBaztF0IHxvrqLEtg/cAeBEbxv3JjTJeLvw7PB+68rLqO9HhJOsp
ttzxfHxpQ/lNgY30WdHwpzaLRd5jq4UEBch1DrP+Kaju8pupGgplCYGGILzyVx0j
BkBukjU2dbVXUHvPNCVGU8FdixxkNtR08m1ze0AYZzBHRZuxiy8iIcYtNKU3r86R
s61zUDLrb3ceuKEwrelznxo3aBYEJhnbX8bhsLQgD/1PuiBV/Qwt4zC7BP8Tlwvp
dTkWpjYReDjny/ljIfA2grpc5W+NjZezjnCjAfk5jQKLOLqAARFB7LFqH/ViSOBV
WvrKEEC8uzkd/eOZjxJ+FctqdKFY0itraKEhNw7nYfJz+hDMaF38y01v3Bc+rRpy
mOVIq0LKztRiOysS7x+ts+t1rI7R+l2BGu+cXdX4rU5ITRt1fxpgp0iw+WgPwS5E
OG/k7uAB6lu8GCfaZ6RBKleSZJVOxdz4AB1zQgH+dMw01gINWHlouuNZAcL4RIT3
tVyq8Xdb54dY8XlModZw+w2ifP+c6tb5nI4wvcLIfg81tt9f11Eoglqi68YRLbLw
2h2F7bpQwNjmjYA99+Jp2WlNf2heC7DSOiows3MPqaob66w87kRXOuvGn3+gOGkq
uC2st2lrhJDOiVwvxhpRAU4bRMZ2B8qhxc6n1OawHbMKaBtKdrLeK26V35hZNEfr
C2Qy3wi5W3wtyjamc91JD5ER4AU7uJ9XTs3g8f2hfZjdRxoZT5bSP1CyfT67VpJP
7fKfULDiKZ4GqB/Qc+N2bAhSPZRT1dqbcI2GXGy/lmpirJvv6fKwu3fgMq55nvra
gXQkCTUPt4y6epSsyMNmXHo59eYF7WoaG5Icw4JonwHkddXlfQ33ISPcP6P9hU5e
KCNCEp6IP4/cDYq5MPXCMNEqdfwNqy9bMdYsjXjtetfRGv/Fd8+eMHtc6Xq+fBzx
ooJd6OVOIhSpMVFwhUd3yvKnlp3B4wfRMurxXSPL7QHBRZGbkSeXdFKXhfhP1q6/
h9ojbCBvkdjDMm1tkucdGejcmOuTeL4Gonsrn11NE/jxXWIPKWp/LBmvQsaZluFh
Lc4S75R6okF2Ch02vFoslfwAxT6b6aZY/RTuFbPHOnQ0r1f/rmwWIdFx+FVqOWdr
OSYo4ciILNMcURIUAIfMiyy+E7yaReXQWpZVj13MG1OHZcAR3R6DGRTb0H09IIQt
QbaVXpN3rYCabUi5cCyh3WJigN6k8zDkq8XA7RRJWsm/IapnImqp0ZHvQXSB1lJf
gwkMPwEu2m6afRGQYHmSRdtpGVVrMETz9hCBaVXNxp/eo5Q4zaftYDquIKznymii
bHw3DdoCwW7HVmD1kgjMAMreNtyi3E9owWOnuWwtrEBX8ISO+Dki7BLCAEabPxVV
DzrRHRff9wG1j/ql+TaV0z12ZtCJWO1Fz7D5HCeyRzhyjykpWUXcFdBSmgpMuwwr
I+sLjfK/ZEfcHhbZrGZUtkqWH4rUTBIqhHvbmZC31bhZqu8JqlDwRi4llDAkuNT5
s78ZFnS1FPTbX/yjK914kwkzTn4uRz2fYj54dDckzXe7UioxZkYxtpRJ+sg8Ob7t
IymjTaZdjldQ0JKChm4nIpndvDTF+XvEokGCEuMTj+oqq/AR4cNtNyhQKtkEIXYS
kNQqsca/+T0Q1DZkN/y7AzcFngeyQyITAlkJmSjLHeCI+JK8rV+lggUbArSI6Khh
4ZhjziSmZfwTqpOiV/6GuOKlpInmfm7+CrcwPiQbMCGt4Bb2l0RRiKoiODbftnJZ
5lKyvvurUuCTUi3q0hx0jZslytJQhwfhaKBzl9gxcZ41JlNYL7Z1huagPgvelOre
oCPgG/xcaP/zmwFyd9bvCH4Cz7mQuc4OQdFTD3Wz0W+I/HPFc/tvvhR7HwH2N63i
5p7LT3ZlXjPOP6yIZn8WXPeC2iIwheNCrVIczKsUmEIk7W6V8XKpDI/E9xDkGoZl
k/C3MV2TOf2H3pzxy/dc1lKUtOowBSSb5QPwwxR02BuR04jTYy3uO3mjYkAXwl7m
/Lahjbx3uLBBk3XaWeB+HoxJKUjrFMxKgGcfNmzDK9Xm/zch8vDhAJA8NCYU2Hqs
B6bu7cw+tN6rwO1Ls1JFx3THAcsIuOD/sO3pJSTxfS8eMBoVTSCQh7EwCYFlnDvC
+JWbxoEbLa/IN5s8VPwzhg0u/Osv+HbQgqEf00wwiSuNui0cuwAk0QH8W0SWMVaU
60F11MjuMN+SeItNu5czhZreqRRyMBisOoQucr9BAoXCnmoYLjWokydrINyq85yN
c85VqKKRT5W16o01oH6P5fLLKnFRq8lKRx14+oeKpfgRaVeY2jkMtpcWIBak8gzY
Fvi41yShngvD0KBsz8r30v7pLEOXhHSR3ZwUHzeFItAqUPlUDk14sauqEYgJViJC
9HcE1P81avQOytJJfqCPmlSDXdmrRDq378ZVO93dXtHKHCUb3M5HQcNjsfxdkCKm
0DIBzUZO9gL/G/IEG4Rivnm2XT4Eh0rgtNe07ruv3jZMIdUwUo1kGKcDZe2NXeIX
M7wUzJ6tXRnDKreJYSYvTwym2nQ9T7EHzGh3Ue/oQQIo4337I//PCPMUefjBsk64
xm6U16Ohzr4ArHImZnmHIKutoq8phM02kOuli4J/cXQ5EjxJ7/w+dD8RR1YOlqeH
RuhgQhY8wW2S3bXTunVwLHdt4xokQQzUK+4L/K0fzWjlto0LvGKJpquBeM13b0ye
ubJCnzEnW68QUmLenZV6Iy2lruTrDmheSTcoiLnhAdCUi5+MDG88ZjevyVzLFQ91
z8roHRkmqdyENhxFsqcakuGeLWBI/V3FrTJ4MLbUOBZff2JQBRaNbF4BAMl5BPrH
Xf7WTVSRAWyKtUhFtmHFI35yL/kaN921Aiu0izPxzZ8eeJ3ILbA+/uS14zzxaAxL
oWzLDjpES0aJd78wesgpfr7fEmoI9gpc5wPE4hqkcCWczBOEh9hKepPUct621NC+
QoOz67hIKIBZifrYDPyGrktzalwq+kyF7PDMrzDZBK+7Vm4xrGoarvMXwtSU6ERb
yRY3oFmOZZR/m3b/g6+C9kzl4T+im7xlXPy7EiH2APXlR9YEZhH1Y9LM1gXaVhG1
c3O98uDr9rnwGDTByB77XZZY/XiYZ2nwIq5JC7myF3rPrS8uieaRJi8M6jS+2VfV
qiMmLRqim3nBNMGow78J73d2UNbeBBNqKzrcnAhhgOGV7AlOU5tnUolTCfVzMra3
2uh/39TwBAZGPAsalnVg6AucZBYRyTa8PzsijiHlksGEW8+GOhinK32St+pNPTah
ZB8HCxB8U52ub0LS+4C8ohHXDAnSh3sNw54e4R3kNlSfMgcOno+okQkLp/ooX1wV
kfQZ35wYYY/jbsAY7zBGQ0GkWQgYtz/Aa1OlYHdQEMR0d5VsxlQ6pnniNCH48YIi
ksbf5fpsqXEJ/JfGIAonM5HAjCe4gi5UhcpXGhEteh1/QcCiwJDORyZdjiebH56m
k08cSC2fFIRQ2Y8YVtFa49IzYNXVSPAHvy+351cYSExQ94DK7xjrlf+QEQXg14XA
puuKybRnSg9Jz3+Vz8AuaWfGjo+ou10D0Mc7Et3xxvOTdZAJWjmH+w2LKhWmp8p7
BYXg/twEeHvFuYNie+npV5Ch0pylfJuT6sbN71UN6MX++pnrA2wJeEn6IJMoCl0j
0FOHf9TkH5NSCExoiYwTPTB9svXZlYxAiHlSfBURUatJvjoox/NpBs5rLONua4H9
Dq5OZQZP32qNezzoztTDSnqpR4oae1rINAzdnjiHbqnj+zyw14qxo0/+G/qGBYya
OtM7nWywXpLJ9lcW+IP8tFmsM+jUnRBNkpdlpN0OsXkxClSjGZyZFLf30aK62EEx
JCAbq20EJcDhivt74aaeBBQE5u0JIDgCnNi+5MOhfp7G1XnkGc41b8YnhYt21ec3
DyfXKS5QU6mDSMMdbmJkEMx5fMOGVmQPdzB9tq+iqEm4L+4SsvcmkD/kg8yZ8RnD
nhlbs7XaogKG9lQ8G7bm/zOEIZ6NC1MWMaElkh+iPQggdySgqkvojtjPSmqCyBxR
O3PGIZU+XatbuCaZ0esDAmeYXqBdJMJ6ecYwxoswxr6rYS4OToUL3qRRoymx7lWc
j0P6lkmWePfI4D3cf+1V1y0JOcmJ+TSmiMLKjQTlQYK27O10gOLl0AXpluX7R4So
njZAg/j1hHC5YSbyZLAoS8rpVhAICRzguOvKMo0jjqvzsF681c4sbTKwC0zyJn79
gHDoYyjWtrl1kIadhhBvwXnwc+m1J7klKyc85laC93JX2NfQMWTGqzw5BOZXlJgp
mzF3xVyW2zQicGJKnBXy8Gy4oPy/7pDsjhOPg43iKWjYC6iSG9WaGyB09Vfu+F8Q
6DwT1yKuBkdNmiM7sGLG01DXsSylR1zljql9mRbU8M7uCdRTPOt2q9zuKW61hU+M
2ZLpIkeMgvRV6m4mXwiydh2XT1Ng8CkaouSWFhRqB7N+PRsb29H41c4gEN+mLk5L
69totQ/JHDPo/b8jP8vY9j2cICntFbfX+15lj7oekde3A1ZMW9XoHTuk09E8GfIb
MuTLrCqouwb+XivEcRObAEkljLTURVZUyLUfj3V/AP7C2OU88gNpPIKssIthxp2J
yhn+10oeb0x341+X5hAz9T4CX2fDEwm1h3yXAj7T8LbgRXcqPvuT5fyH9QJKWIOn
gUF+mO7thrdj5gouh6ffzTeot2U6xCSeflzY/TyTp9oOEYqOlB5Ck4AIVx8IJSRx
KwufMevnASliFXA0dKzfZ9OXBWv9cwPX2tx1ALAsea66EsnoTanw1lf2mV4MOVCU
aizxgQtP7a7N5Rw5T7Re8j0ZFagQSCJqp16k71XhUnroqSG/G8wwqswW3irjV9K3
NKernwq8kBbFDl/O+6FDablSpehHLPPee8TYxvc/vQqCgEvH2nZR7OKKcXReDtEp
0OGgCWGrnAITxZhnsMgE+XpqudNxfKFWtfTGxMZ19S98HpfbeSV9FatzwboENsC0
DtcEf7USLUVTXjOKiZfwyYfaGrIk688RrhlOebDx5btFbMGhCKy0k6a1pHrzm/kf
e/DyZ68l94ZVlTwEmrMvLGW2oh2asoaz+Tzkvdi7qNwFRH1tPE5hraz89y/ESuJi
LHyWcWr5NwAqsCZdcLCRNUWjDPw/vrHj+0/QbUC2mo0+Ky8ROnnraPQqyqm+5Ck2
exgI03BYBBz1jcyv+IfF+WHuSRlqxpZTbgU2ZCSdoiQwnvpLgd5k3OxxgESjRDbz
JooYCeQeOJib1ux+xf/v1tA43Qe5n2BfTgHySyLbiDGYjSJIXakyMi3xqpr/pKjc
xiFyAJPiRrtpBdx34DrcItp82PVEWloE91z/NJBGtsGKOKo2LefAv9s1q9IaEL/n
WdKPEZ4kJzaHIitL09Ev9RVdJrC3NLUixJkv31b/TaxPnp+SIdvIkKdjqZ3T2eT7
E3M28jkYyhpAqK2KGd28+jqRGQlB57jbZHr+ib0UDDFetWKh3QTxCgl78sahRIvw
7NGrtc6x3sw3DTC9I9/PWydYlYc+QzBpydQk1XkYS5mwISChQzvMvKgAORtzQVHs
dn+QhhwE6SBeoQ4Tj+AZ/XTQNVp8NIIBuuhoNVCDksfC/sVNO+5lSj/fqAhXo5Mh
Tc1hECRGTJnI5byJF4vgth84fqb3GJZ54zo2fbtz57/VRwsPz3JM4HqozsYMPUgh
6CgcjfhmSa04esj4Yr2WH0aKVY/tOQQyuUR5aBfxSrxmMybsSVzcCl8KldP3D5rT
x1zNkor89vp3H2beFeSWDnaV4Y0YXvlfnP8/FHJD8anDnOmyObOcsApOffMlp+ih
dCVqvEjP2+LyaY0fLCBfa/RYCS51BLPYUeklNmHK3FREdQM4FSf5qlsTz0NEl+eq
hVgAXkhAiBEO+3KGgRwBbZLDfjVaQycUx+wki7xa3yUYYvkNQJdGSibNGll1ijLV
dxVn7i7wVQeHWhjhk2oJRqtH7dhEb/6VqpZBj8oMob9P1QfF40h0oGJCoM/3BKD1
3iOym7/sAlf0VcCUAhAsuNyaybySICorH2TQ61YMYBa2Gp53kg25vdm3MOU0o3nz
7P4IPGcSqUSTq7i6gnHJY9ugWFTVStiN9inBE93e6Yp+5KCKbbOx8oXNvbWHFAb+
QHiDo3frLbu65lS8+nU2hbQGny7vRllgagFaYDhWx7uereGOPiIu8hJYx5cQZXhN
OvHUM73dkoRlC1J8GZyB7Xy9qqTvY+hJx19K8HWc6e95G2lXEY2GHub38HbYYqH4
lLtjorjeUSdKX2x6bfy15GN0hn1e5j5rKrpv/TjX/D4sBbD0Mt5/pSRz1rMZWqs/
xrNPNsqiRfxrRqdGMTvwAoWvFxy1SoWJR4e+t2gT+qIYb3k3k9gCrTl3hiUy5A8/
bTN0xO4JhQmLArvUx8Pe1fsuGYr0Y0D1ECqN+gyF3vZelNnRyiRHuGSB88Yxzq0E
jbQ/5sQ42QGVuSWXAmiCAIdLuDfWlo8R8kMx1xaV35eQJkxIZ0CIgmfJcMDH/BMv
VdsVUsp4iuhW7chaWr5HKWpA/h2FhOZR4PFg3Is5jGfnjLaLlxMj2c+93LJtQ/el
6iXBpFaJ/qyDlh3+7wOPVTky/yOBYBcGd7++gkkkhAWMxqPCe4o4X21maJvviZ4I
08rXWmFvqTF9JiU89OC4w/kxFUojuMMBsLu761SeBb9ub+ZQn3B/fZgfQjT5uyQu
hl8l0TYRtwx+f4QGip5lrZF2TSqKbzCuWsas1Le2b45Dgio8jhKAoejFnIxWiaqc
VuhGL+KDUpe3XPIA3q/UnU3kXtHRkOEl7FZUQNkBKPLFd64QmzH/ySQw/dtdIiUV
Zk6NJOHWI44S5KI8H9TO5SPaESJAFNNfYAi5+QOyZmpAkhzMLssnviJoCetG4w7S
J9e1Mks5OEkl0uCEMwY3NFIsvPkHXVBYZqQyHiExAcb3nixQ6XfpmJFhwf+kZRqq
A7dl9/PlE/Q17UgsDfVhQljnB4tJl+95O00a4WDtmO0H1CtSZIKmAG+S+L7o5OSQ
8IjUX6t7e34OAyg3HXd4RSxl4hkKRUAnI6ftmFl6oepPZVBxsILfmze0kqo/MNRh
ofdx5hihYTaZ8cYTG9fLTZ5H25ROW2HqddzQDgx5zm1cFwvT9nI9U0FRrxosqNNL
R2iPW9mrT6hM5c5poV9fvB1znSgNtPGitfqbm/tzFRMLOnhJcw4olh5kRgRNCXTl
AhAWnlJCG1rXTWTMHMBtKu8lpIAvNgr0mDHaCN2zjIxFKJeqhA8HebVWfsBI2bWy
MoclpWdDtsV+Zxlfo3ZAsHU4bsVZvELY2pFgK33prU+nKK9Jwpb+/qOmhl9z+GDW
Qhm1P/Mm4kaBQ2XCiazG5OQttDdZq/IsGvyBFdEJ25o0dkbDwaUXS4wC2X7H/jRU
1m7kV6/STj2OYThF5hTi0qy/RoZJnChgF0+guPTPgcZ6sog7G6Kcm9FGk8mevRle
/kLmxlo+Ux6voYDlKDsWovqD9Xy/5sqdhxsaTqlhua7sBLx+nYlT5O2qxVY5HAuj
iHjwO/nVmLHhzzNTkvO3izOx6id6K3QN7NSxIZGkHpmXA6bi8rNECSBpLgK88aiH
3RcPJvflrdSuGwWbKO9G997DUTgTQpWy3jMYWbGE6o6Vpnjwnn9IYBDMiv80vpMN
/Kyn/oTZCQEhC4lDbmSlhaOrTtPjgP0AYJu4naq57QTf//LAtfW9TmsaYNplaSWS
VEBmD8Nvujj/oWUm5TgafIR/jt13qRD4GRxo7nONyQo1tGUUVkcsBs5ZSOTOAtNw
7a2ekoyGE3OwzPjcMMpbQ2iDBRhNVCXew1SIAAOy9By2so2BRTNpjq8xW4Ciff7T
yry5YiG1oanDWEtBnN4a7C7GMmfyqK6pz1v6r+PKqIXZFhHwLxhRWINJtKEyGf5U
XVDxV4SoCSZLr8HKm5x0xc4Q46p54WeeBdaVZvRb9TDFVVW+bvALuLA6krAPEIo8
W7WZkYcKRKx7kj1/de+Knlkn9MZ16kjVPNfLGGB6sEETj5hfhhdcZVWwkW/+CEvE
H+6sY5wRdeTsarHo/yJQM0WGiFpeA0CmgQiSeIJZ5WWXsDsRY7D2h0doyffyCfWb
UoFyFDRv7vp+wcF9OY8cyRYU1U8iHi0ieNQeJMqYg5ezPgqWclABc9O1jTQwFFLU
5zpHYn7EEKwpuXkT6Wd5z7RKIwEEsa5aItliGxS58wdtP4K4SpT6Xq6PasBwYkkf
Xf2vIV1xgDEkSnjvy67YLdh+tjuB6/mW3YvcJvbWu0konRaTBsLFgZwTOgagMQ1g
Wa4FOxL5c8Z80IJK2UUlrYU9bjkfdEmhvDw3sRrWv1N3+RUUsKg6XKqvL6fEo08o
Afk2vVcZsjHfa+8APLiDfhOjQo9viEOC8TGpR3L5igSsJLLzl1g5sEqGY2aaQ3Is
KcOIWf7pKABt+5jIsX1VlP397zCfBSEz6tRyNCGyWDcZfpQhlsGfna7v+DzMXuoZ
qccxpGKTkpvJwZmeff6/DheTjfTHXIOK24D5Pm159nvXUnmAsvuKs1vnfqF9ScLM
IEPhFb7rKHI1+0r6tleSIYHCar/Ry7Qjc+kZviGAclmWIWZSy2eBWhzkmjB9EXQ2
C3+p36Nqc6oS3Jab4bbibDp1JdcJJyPE4Xgw9w7tR5THjHAyIS/eU+jmpKz/UD50
Sb6BcROOw+wiLB9NvmHnoUz58M2GH5kki/BzmkF5pHfgHNxQWq/rTXRQoG4k9Ecp
mEUDmBLo9sPEdUvvRaGmoCu7Pzveq91Sgz9UQNT4fgQhMuUKTlCC1AtyydgodADj
VH9xGC2aXN6rkvQ37qsTbTr95ST+d4JmNMHe151e9BJvXuFGnC+dY11jZ7KVneZg
bkye+Aq7th/8cczcKjjc9L/c2ycpV6DF4zNzkiGHKHoY72/u17bchgzbDbRiLcPz
XwIe8E52h1+d4RIoU+WZLrZs5m8Ol+POrNPydhlEHIQG3xduKXc9YkVtOxReCJov
wNxxMfBku64cPVrqLAQIc2NV1M375DpbQqzfT53gafAZ3hr8Rnu1ZEQJPnCrtkdX
y18Pnsf3IxLi34ODl0KjpV8cIsPf1+qVLDsMVHmQ4IgU82UkQsUSZiO7Col8jqi7
2hAa5QlUb0Zzl/NlGrIYFsXWPr8MNTzLHflmTNMeXsyOals02rL8dueanzholoDl
TpyYfmkNRQUoYcUZYH0+xiGCxGODaWrCOwEsdb0RQdK3HQwgLycO3UNxgYe1K8pa
/xfghIJgwvtu4Fbpfa0CPDP18kLo+sfHjYtk+7Gm+nAg5kNrfG67XPj2DF+v0iVg
nTc0vnrXhWdPTfPNUAPiL6Jq1BR7bgmqI02QPfdQZfOnwOEVf7iqGvki0WFZCd+Y
74LUcrhPW9AETep2tTAWi+gcG829d9L7husbtMDTc2QUhiCEIwrhMTTRlz8R9FKZ
N8Vlt2xTZLzcN1Y03C4BCdqHJjB5u4uz2PALKoge0ej+0bEklUhXbHXXSG1bg5NO
c9BY3FFjXbCb+bBk2jTzGbJXCwXyGFN56X+mTIIa2GoVVs6AtVoUBB+Fr+I1Rrnb
UxThWKgbWau5W0GIxzEJwVwm5Gdr6/sMhorxhu+QTvB7/0DWz0GTg2bdERkys8gC
frzJip9AnMQQpQ6p8LK2Y379oZ/ZdcH2FVYJb/ZigXR8qYegD2UkiNSaQUDhrLS9
7n2yHlrDUYy/V00aCTA2TNyyoYZYt3N8ys8KxPcH23BzsIFeWTSLHhbEOPHrMnsw
zobEk493FrJ2FY+r8CvE7H78DpzDvxP0VAzPtdLvEBO3mAjXfBmg/FR6e38WWUzj
j+HiN79+v+6P73n6feXb1bMYt5m7ltBV2Hu6Vm3aoZtF0YXwhO8lRzZl9gaaZ8ii
olq2IRPktPp0T2m2Aw4WubmJPuBX+ITGFubs8gteXtvtojZZiIafwgBp/N4M8Omp
czevfpC51YLD2UvZ3DLNJLNJkzmDifLjaDtXt9eXM0699XA/0WgkFcQEmfIk84Qg
89/VZQGQUAYNpq72+vMsMYhoad4wDplZHobJFfIp8hA838rCv1ZXjZW1W7NBhicc
gFXF7j/wgzZMc0NHELmjNgLCMRLkN/vrecB69MWHc5CsOXflvxFvQvsr6Gx2rxeq
3Njxc9pRn4iC8dqSrZNOE3gsvP9KmwOprzAKPxrCVGu4Ylip5jdTrsuSISp/tDQ/
Nf7LTXRQHnML2EsplRw9+O/E/lUKT6zFVWwd8zHoQfD3rX9/Ez8KOq+LJ+mwjnSC
RQBXgG16X2rmETfEieLPbMB9iH36Ai0VuQLaskXTGEjNnR36p1sN1pmlxZr+ogIn
r++mR3zUf1s3DPW2KBt83SirQrg278IXhbSYSeagpgl2tG4JRzGoLePAb8E+49AY
gEOzzWl3qTy7zaPwvHdx8yK0JrS5Ncw1dC5bobeYB6T9/ERMoYUE/80WbOWnW283
4wLJ6hijoykusS3VGzkRWY21rMmtPxeyor9RYOTh3971VBlg66LGywnuJvIzZLJh
Ok/8aPkTLcidMYvTHcgQV88yRhtdODZfe2xWLOovdOfWpfqIU5yWC4/R9iphddoE
At1EEeQckbtjjG1MurrA/Lbxbn+Uqv5fkF6ZwYGKsOhsolzZUvD2vVHnvIZvWaSu
P7kOOthn0BhpyMeRYYlo2Na0byeZVaspmxABM2Teb0BXFLb6UBydjZs/jZQABH9l
FGLF2W03TW8oUfNG5xOLtyGnWfeZUZPcn3CLawD0wo7y6cismTpo+ZOlhKe5Kx03
c/HDisgvLoiG4GsfVlqNwPB844omf6qHSMTNwP8Tx/xC5SWbKyHcosjfGrCO9EC8
4XBk2ddm0ScVBPEeV/iy7vwBFouKsFcRyz+ck6nSIi+C540EuGK4XjpcxiLp7rZj
GTYQ1MWZoZ73iyaf8Rp8EY84+b8oqpDC8tV40DM4rWoU8EYVgoF+at4UfmNMhhOJ
ElCV4IovD3SZ4oOpJsN77bh3e+QuIOEXHH9bB70sXxxfw97w4KYOHEUIXxcaHe83
tnMXDK0DCPBBn6Rjivf+cDGqKFy1iOknelcOWSaPsbC8fLiSJfaX2tAbo3FjoFFr
5cdUNw93mdv0Pawko32winO68PUKrM8AjueeCBQaLpBfRYLxJ0twzj1sz7rGKlUK
0gjCoATX9AmX2cwy2ngeqX20ooPI8VaoyGKSd7gbGqURhqDQxNODkmQH6mympNS3
cCwGMMiIZ1PUgsDRk0RX8LazioQTr0Y8MCVYpDHaGxXQQaJXxRQRp5kCWMwK4dla
83pp49XbEZTNzay01Iz5ywnKcH4UeAMX7SQA9H5r2kTHw1nsbG9FzB6UzFvlstvG
Ja70AtttFsf2uCxloDJeFpC9lr9j0jTHu5bDgbtaz3vuRou7XTpyLd4TsgwGWclK
kDfMLYVdVXyEkJ61aw2UnX3vugKtiiQu0Wa62uZC0nVCHufU3Nh1+tkSHdh9Sbis
B7lOe6FNc/TxZgSV8fQFj6T7Y1Xwi/NkcCC+oos7ANHhL43wLCcQVJ9NgFZbYLiD
DRSNuqt1kEKHOp4HxPTbZRscT4X8bPtEaCRwV7BjTd2Dpk6fgBWyOxzPz0Vjn9Kh
H0gLaaQl76In3gwI4tmPh15Y46r6rwOrSkFk8YyYu19DHcrfCOXuZ8FrUJRRhr0U
VKgFoejhfUN+EvF2oBFRaG55JKfl5aPDCbc9CAJCNP73IRnnmV8QWmvLj7G1rcER
B3dYGh2Di7AnTsy3mL2eGKnrkhsGsneyQRuObFNt8WCUQ7jhKoBS9EPEXRcvSMJz
aOWFs+874c2kBoQwAFiXFDGT3c0vJY909srtgTPfWjRyF244wQPKd8rjYbXgUb8Q
QmKD/KHh9pL5nPb0PTwWJdtiwb+8DcXitgrt72ksgsa+2/JqgtC3QKYkjre6OSyU
S3Kea2tU2KL3PQSkQAMPUWwHxLR+fvA/RYzjCzYzRmh80h/UabggoONUF4je0DD2
rAAca050rKRzbJPB713NH9sTnKxxmD8nBAc56c3HxWhxaVitajf5zAPuiDav6eOn
/maN17qLkU81lIf60lNlJld7S4khygP/oTDQ9uyDNczzFn0mstsTpd1yniZuPHOT
gSGbvWiHUoagLuFX6rvMaQWnKBR8w/hw1xyyuK2RTMDUlQgBC9p9aaq65wrMqBNZ
E4hzFMCFAcSPa+ZkeWQkqktx0EJvKGoUmy1t1rSjlZfxMVIhmcicwQgC111wRlkd
iOl1vf7r9v+ktwGAnwWJh4QxI42HtKUamuHFUZlfO6EOi9x/boc0f/j15ySWZ+Zq
VRbELuofGiOuW2w8XMNcXx3eecrpvVDDiQEjZ1qwkbGrpKeDXNZJkoqdFeHNm2lC
N1Llk0/j30qgSfLrxtuTsBWfjgOHMclYiz24hNavSceWs9Nr4sazlNplLzVURNfr
nvyrUVXHprLUmY+yLhyaTo7DH+OPx2SPzfaroXiiDj2MYtNII7vdq1mDPphjv56R
GBtqs8hCEUkg4PpG3K/ZWTCmvODgQbFMEVN2KDpCts74/4OjuUx2nAGH1IeUThf6
EXVu+ZVWLEdcMQGc3CCRKmqq2/JMr69tn4Hug3uw6al3geT6Nmkju1DyHnMpJAA1
fPMTgHQF80qnx3PhDkErL5oUDePcAdH6dv0jLHJtqZR7GQ34R2u5AUi+/cT3zfCE
/d+76Q7Ur7zvitcZzcRxy87g2PdDc9SfNbUNy3qmRGtkp2gYKxk48EkYoRHv6Zd/
nba37XFHN0bGaFstg3jAczNQ1RWzDIL8NwvLdlXGyt2P6xfWg2tUJd+1lpeK3UDx
oEGVgjRW5ePhQY95s9UHOqScxEFGmlPB98QpP3KfnGBbIA6tk+pFn72KIm0InNAA
9G1GV22oIHOhilDcKqDT8kkL22i5drhlwr0vuaiGoagJ+Pm885u+6l4wIjpyGr3W
lfxVhk9EUoADSZ8HmOKW4Q3muU0xQ8uC2YvB91PQ3WyigxZ9deuAWZr0DwtwkCZq
V9/LAIr+loQ/+s4j6MaejN/27fqXjXJQvnL7WZHOia65cmY/VsxEsn1SCJtTijwK
tSpTteWzZqHcSQ7xKG1hDuHQ/bqskozWynKAIuzd4DNBPXzzBU18vDAt7Xlj8O77
qV7PsTqerdztk1mrXLu0K6WAp+4A08AvkGqZ4m5Wjhm9lpr6Ay4Lya4mE7sYuSWW
+6/I4C3px2m2XEDUj9zTGHsKpwYumYGBs4TCa0fEnRy3DQpPSnRJI/WDNGXPSi06
ng/RHsHjldOJVhJ8U5yWV53Sbn5IHOoYr/Mu78Zb/nc1426nYwhgegehU50YbUTp
+t8XmfeiOoiPrrRxS7l3ODXiMZtpHURHzoIdk6Gb+OD9XwH1Tx+BfTcOTVMe0ihR
oBPQJlppOvAR+Ia0VWakFsHrfWfmkxthx9jKcI2yVv+qrDYxRKqdcQRlMF4aqQky
UKd8SpBFf7M7qMnRKPT9p3w1MtJq7s3fPChva/xhSlpH+cJ+IWcz7NjFQtYqWYzm
4pbA4wog2FpmhVs6Zymi/nzv896+gcgYO7/lW4y9x8zd3gHjuXVFIPgkpKzcA0YZ
nxWjrS8ycT2A8JfevAd428jmNZIhWNM987SRTjPA3HnvvdVAoOwl7HaN6XEh9bsz
/yK3nbwPUpC1X/qLGPfZLL1j037i5I2SHDKotx5mhhOsagr8xu7pyhABYwq6UgwG
Vv/jfQo46ZA1HWQds4kq6Z5SJqAttsWpQ+X+oROFp8KWVsuMvSaxKhHoiMgstbPk
bELMrbbTur0XyVWubYLHJFMOflwTZ3gwd53EH1LMLzrz/bM68fwusM5iSKFQ99YN
6qfsrDVhbzlrQ4lH8oLhtOwzKOp6SQwDEYBMHXbK7rUrOHnSkSUrqGtbFZ5Y5lea
qjjhJuadgdp/yiIVemGgIUdoOvQoZ3p3nJxcIlP7G15zsEPsjIDyPIcGwaPnPoiy
azoODINpDpdd54EL+ICWFr1TUwksHsk6FuQd1YRbpq83gSsjwqJ1104d/7MeTVbD
0XjiOZXZWsEavXj714aAOAwwnX+RUW1gM3aiiCnnN38EF7FGFdWQFE1zzMa7Yjqg
+AucWJeJAXNMJP6BI7snMTVpwIai0FUg72j8ecYlW4B5NrHR3KRclc+BuNYycYwB
VzPFY4N7kFv2pFCWEfX2tHsRfGMzqAa1y/d2PLQlSVos/4nX7CePH9YIFuLMNu8Z
dAfHyTFdJteFPiMVU021UtvyIgj3qlWS2YhaGm7Un88JTFZJ72HsLpn+jrF/beYH
fubiIvpKKswOAnRN6G0k/vmNMNhwuFRiCMFDM2jyLPzuU0hxdl9ODEGPF0z5X1jS
mC1UgtDkPQb+lfKUb/zjP0q7H+75IFcu+u8qPB3cI2v/uJVEVYhWRm6Y9pc3pM54
kWujviaZgISmqGT+VXaKpDKDgrgj81gsqHrtt71WfrM0B5AvJhb+7kK7Vo9wUFwG
9px7KBa/lEcEJdZKwIO1j1u3+k04UvMkUsLhjy546E8tNWlOClvCnRtg5pV7mcpA
w6GBIa/CcrCrGgkDVnLItjsD193/u8PgzcSgDEFpuxZiWJsOGEclaSYDI8UfO6m/
N5JeKMvI0WyFtlFbGVG3a0KZzsyEl7jU3gjlHbIDi2r5bL7JJ5l0Xq9kH0zBPgYS
Wk4kv8t+xFmUJSL4oL+J/5i0jQFL8Enmz6S0yNRM9fIXoj+qpXfjmghYBfHCF5kM
Owtz/nplHW5RXRC7dPUqA80n43XeZYiAB+gTQ3il/Fj6rgUCW6FtnLV5++QuJnYh
FwW5+ZVmqaiu556x9mOSvrYPxUfdg8PCAXmA7GzdkUB/Kz1Pj0saYSmw6YvODLpz
cB7vkzvx1DJReYE0iDaMlH3AKPmQYb5vM5nZRiFqIJr3k5aGP6RffoD2JRrZF4x0
fZFy3rtb9Da2fI4jMKe8DJ8QBWGxhnFk41kRN78FhUozYR5zQWOkrfbmneKBxT9Y
TdQydOMGoSCzFH9NhxXNnsAclBy5wjHWCU202aaNQiNr1bSUofZAwBvsJcmIVXVL
XNUll3CTaPDIgVEXzoViYyFdIjHxK+8XC52LVeQKc650jnthfcEJ+GQNKNP3iYhS
l0rV/0rNkzDayDU2GFG9KBjzyoGmvuoylKgFWekWNqBP21cTspD9+1iPQgoEFr06
YPYK3msfjCTy6Bpou1JL9hRqQP5tZZxF44SQhiIEAZserwm+xTQ3B/Aq/RNkYldp
bi6Uui8kUTk8tuEyNWWdlNs7WhAPPxduqhn23CgPZS/oAcF9AcfGsEjYl/hrVC9u
CIZbnQSBz6Hfwb3QpEQWk2SkxUD3GPv0fWSnOu5Ri26djwvvhwfm95MgGGbBdw0h
HqnSL7YIlVcBISqc7fdudftAGDJhkYA4hpAcUIwORAqFwinAJiBglmPt2poLDV0W
kEkxEtSnszIJrxMtXKhwpbNOfoDiBEWXh7DyPKQFpE0BzgHKRjYm8NpYf/cGA4QE
INBm87M8/p8xmaDdAkalxIHYpQozj5gmyJBPGC9IYNKX38zV1hgNs09vgE4rBVci
cowknQHecapmsM4jLu128v3cgrnd7Wfqbagmq5V1zhNHotgXGs+/TOef5cJCRUrf
UwuLJdgqqMVkCuuCp27XQ35G7zsFONe02tySCM2QFLTw3aptQ3shmvUqQRMvA+mr
WrpHome0OFHzjwXY0NfYfBVXLscYLGbGQjw3dWnzjJniQuDClzoE2TFtP3ynH8NI
1D3B8MlxAbjXkzENZNcxn2C7zMy/TFlKxuJ7xL5Ke/jtBD7EGkAGML3V77gd/GZe
Mb0OQC/9iwc8TCctfd+4PAZSjY1KxvMrL3cupEcrfHM2WgS3l/u5NLG7q9m1gcON
gWcXOHO/4/zVwImn+5uX8Cy6Yt+dKiWA6O/pizuAnJiq2Y6mw7Ps1vOsm/w3BN95
avLkuD0RfDAXQBnLPBYQEtdeLrmDxhLIAMW528wbPBbSqF6e6ZDF9CZkPoOWXkrR
UZ1yjM0m42xpAJxzDPLdhbP7Jom2BvYtsrAe1i1qWdpnPRmBsDprowntVAMuzVUr
IBvmMZFFylOTdCUnf/etMMkMGPxv2Eb1YNgjbCvJsIDMXTt36n3/Xte68w5TUtUR
rRc4WmHbCHhQG7qSknFvCqaGQirj27J5AlZiY3igAo94uIgPf3KKTtM7WgkHdX5w
ipdU5UcTCrOxfqfpGlLn9ILw05usO2V4HZal5qyvZmwHgXnHy8/G409L3MJCEbVl
tqDd6iEIKohNXxp07JWlr8ep+V9Y6grTFTzRSF7/DPGiaKW4fgoJTKqq644OcjNo
NuEHn94BvZmiC+k69guIH1W0NsIEkyyygVDXzibVLwUDXGAvc/nKj8gAEJTWi/fK
8p3R470aFHJDURNGWUjTMTeLcxSr7i4EBPR2Cs7Ot0Y4r/WC9xwMDc626ux14ed1
O+uT3PZvFmqidJYDDIk06A7oHqt8bUniN4qLlw78Z273XzoUSY42wsAvyBhHFQbL
gLZ/H1Yx6Pbj4BwfpyhBHHqkNsiT22mf47MhEtX5/epCfRP/nZ1DCtxaQZ9H7lHF
t15H1/YuvnE70JJQMrUet0YUpUIGkgDR7hTdt6Vw8s6OSkzWpU7ZSBc3FEDAxtGE
ezbafW761uBMpvYmchQzgl0BKRUYkBdmWg9GDR/qqZzLUEC5wOqQwHW6uoqdNOMp
2gZ0t1a4nZ2LnI3wlwMXAMNJMDOxLZ+6oR7mM8scyc0i6vQY4DSLU5a6Hlv93cvt
uvhsRBUsDGJQzlR9lHEMVTGjjonUzye9AiMlI8mgm4kjJITnB0A9G3xVD/RRxfKb
ifhzcLaMepo7U0nXGQwxYdKGlY0dGgo+ftigFC//fzevD9K7a935atPCRNhJp2U+
2bzccGz1GZYJljLdXU8+2oK8PZG5JSVf8lwZZy+l9WMbGGafdPYDwoGWzMj6A1+y
OUrtU+pHTszTr7Z8GI1Z5wUEs+UK+qFOEjPmLoq5RbWVd3CvRq7T1ZLnFvqDQRyM
1MeLTIYHAH7TvpmtuRxJ1YV3Ne58qCcDrP7rsrgWFsJfm5cZH/2/+gZinFzc0M4u
FJ//C6lBkJbqfirOF2oQ96HJSDxbqjFyszGJWPUymCvI+akyOvEBS0IGDIMIrmNT
CYeO+IPVdUtoVpF6xhgr35AgqB/WXDpwbBIB8QNLsHcrcVbIz5bAjE50aJykzku4
ezRdrixzQzMe8wKF93DtpW8uLTTWH3M4g/SiM1Ze4b5xIPN4+1W48MVW1maxJvkV
ZYWGfMoiH4l1qbtzD7cyI+IREiLGP/xy+01hWPLLPAmH1eSH6ed9P0lFLdpoylgu
tpe6jpE7IWmj/6nVBiE16tyupe4tgiRwGQSqA3NCdxT5kChi5+h1bL80gXRds/E8
JkEMK3/6LhVJBLW1Is07S4x/saFeeuBk/yLid/XSy3Y2c46c8iGqNB8B/XfPwtrs
UbpTK8AMzggml/cCe034e6lP4MHdV872NcVWS4NLLycFxTUiXxNWRmYCf3ZHHoaC
FHswULl4YvRzIhEZzKpruWIfrKibA7Pun0xC0kHwSkH7gXnyIZo0v8HtXDoBBq9G
iYrN/YAhU2JDvfOsGtQ90xXSWhe654vPZjET/++/fLgrt3K0Gc5fk779VPehB2IB
gvlhHT66FNzBmv3DyzxsTYHk1rRBKf3pwMqusfzTY6cOKZsRFpAwDLGWpBP7QvYu
zel8DSNZEzMh9Flmak2Bth3VQMe5qNEusJUbaKRWjT9mIi7szdiKqqxMCnnIYeZ+
gPj75GrD0pl5KURm+4L5mtcEdZJgrFgvTiRUFWXCBkXIFpAYpl7QSflDb4KjcW6r
ZZqmhnBVC2cIKUIywr78emBYkMj/qDY4NgD9yEuU8KsyW+5U3NvDzDtg99X9M7wH
t/Y4KLpsml3b1/G6QzoZkZRc6PWnySrFnXspl7b+h6/4QwHx4bnVmNkPp54HGc/V
oQVEtVzzHuqMfFKcHQf5wBKkwZAH/OSWadehpr1Iz654Tfq35SEFJ7TV1DWNQBXr
z/MTgjrwzNqoKLRpLp8dJI7kRvs9W+YKJGzb0Vv8PNufIG8g8QNTMEmf3RH4O3jL
Vub1U1EmFrlYZlcASsK7/wlhisHiUcSb9YVsj1LR6HnVK/z2D8VjXKS0Uz3+kMZG
m2AIDN4a/KO+jnMkLpFIQmvlyZ5qIU39UfYsdzo3g4NRAbYNrv+oPfQqifunfXyD
ECoDRZ8ZBcshau4iYDZMLgyoriURZ+GXFf261S0QDvVAD5xvwZO3G6Xs7GvSzb0M
HVTJhOrD6JtCxSoUOJQk12kV4acQca0rTfasAvtjlKT1lTPNd0KS4Vu2aD4YBzOm
wK+e8Jpdbsvd8+Ovz5X74BguNXaYWl+C51xvA/3w4rRApBDO4aMpRJIegtg1sZR5
2IgNSQItVbWsp/zrQOubvtW0tiYQr2jRm4iWAQGQ/QGiH//xL5YwzVKwQ9tElzDg
/Xu/cGrYhP8PbfgGlrxW5XNWRt7X9dDzNT2rxNmPuFAPgvAA7Jgai9Q4nX1DfOXG
AJwF4+VW+Y3xb8c97ag/mspSqhDJTecmXOfR4eJePmIKaryo27tyQV6EzDi2hiXz
1hUCU3n38ekt0ZF3+75FieS9TUQaynwsqMnzovHLRDp6cqQXQTIXb9FCTHiZTmjf
BklW89Za0rpPm2LFswCmpt0a0EKUs+riSdS26RYgtzqBw4tNaxhywSyOQ9b082j1
iDXZnIOeZAgRrD86OaZynlEG//vwKs6KKIM2s6CRWd01UVCO2oQ6KIUd545+E53b
oxlAA3i6z/F7qPs3xInLb6sOQwke5MMlG8rV78Jw8yD0uP5PmI334vZ+YkC5VwYq
68d6H8NU34vxlUK6+iG7vbC8hXhNLoYtUfs0+1d01M8DPfGnJ22FWrEIy9Ufv0y/
l7O9vdYmuplKC3g56d8obieIW8q1uyvuk1ZuHU09KgcryLsCKRPJs9DKw9+HFjPa
70Cy38CQTWYrG5tfEyPfrkx6e9BLUhvyIKkU0vR5OQ6q9+M1dLndQq7VXRR31Gud
KKTZXumOx8xvamSrbCeQLy6uuWvI/znHBG1Em92/6+oWWk1bqiwxt8ss/S4+clCy
od7/1FVAmiHcO+VhRdEAHsdeQko5J/Bx+MXOMaFIrZ/+838me/4XG1bXHo4etaFH
BgoMWBY10UwPx3OKhvztkbb8HGXVFV+5Ib/fsZhcfxg5yOQJJaNKvI89XdVjoVA4
7q/wef3bh9FH8pmzwiYTEYK6EWljHceECIBjE2Xj7ou8AqMKEnaGvPSxgjkeIWg/
shcD5q6GvAEAo3KtDeWCGGs4n1zXQI19+/p97sB6vqKO8eOnL7Rv+uX7dcmGLfou
RTKN9Ly2RlsdCmmO+JtSJ2zh2NZebweyHG6IdPKz44mardOnUKcfztetdTDuTPYx
KQfnyf42mvs12kLy4pKZMnFcod/kZQz04dtwNDODEF6e4lfvJ+9j2cvvC/rCOFV/
q1ZHrD1B9tw7/1WQEpcEsxG4yrLK/qlt/FGfpyGrWHGhdaTEbSnsU0y3gxTtw0Hf
H2j8petk4ZeqwUO7QWYeT2xHtzf5F+eiBs27MNn4DJrhdZCgOhMu8zftu+o8ZHpl
0z6wG5DCNp15YgZzov+oNdTxyXiT29P0Ecw8uqn1HdV198qMug8DJBVXbJMjQty2
8EnlKvfbinpgvw8M/iUkxTY0A6e52jyJfoEhsn45XZBGJ4B44JJUBo/phJiGU9ap
jSIo7MqBa0bfHCPwJ82iecQXa5Vdtx14nYJrekyqaSnYVd24RYlCQqObqP3c0a94
GS+vspztExQyUC11qb4ByHSxqyMMeZnrjYQcFpBVWm3D95Uqyoqfua4B+Plr4fbW
KAMujoQKif7iZa/pVCCpSAj+zoDFfjzFjXkLmORxKWDShK2oqT87IS3dR5kzWRWe
ZVoJr82ftPdzw/a+5zP3y0KmLlYMrR6bNs18plPiRUoHYXLz+QQXqWfnnL1IukKG
5mITa+XXi9+Hc3TlNI9+qODXTR7xv3hZG3pJr1LU3221dN9cwt7FOJz95v8wJpsj
C+to2YNajitP3ACPSOljs6C+wBylzZYmPo4fvaHR2AFl8ryzNCKUZKLhot4pUyS/
fIAXvHZv3aNAIQAlC3JlUw3momwh33xIWsyAmDjwElJrqdMT+XxFDsIpMkBIifSN
Ugtpd/TW4FizcXo5BArg5lkqvbZGb7Jg/s5ihkXYYPwAwq1yaAnvJieekaBQ89h8
R1vf1RLudzva5RoD4/AuNIyibClX0z4kSfP8M+z5YPC4bDuzCZ1DRS0Z4mabL1/W
jbkJD+XSQEXNXf+OIEuUpGUKmjYPPWHmMdgVZLGUPOk+W/Qw/o+zP3aFqh+3q3M+
IUPf9ZcDiniXTX3wuKKjnt8nhi4bOX5FXJSpYttB0oS1QkosvZDId6E2nq1ZUVPJ
U+TCd2JfVsSomXHdka4OIGv8JRoDRTAyI4fPrinosVimenZNM7aPB+UlVqkrJ0Nl
h597ATUjbhSdgYDawRkSmfNWqgbHsyZHE9jfXPyHjUgxxnuUtFoNz7p1F8I2uxpd
hhW4dVSERYf5O+xg2E0XNY6FE4mC5IhGqMq/Qcuk1UPd5sdipla7XUNcUg9s4aeX
6TWr7NSUDoAlWNHq5R0cMiSrVpcliB79oPe/hd6Wa7KDXY68n5wx/V33JSqQJIuY
2V0Iy96JiEMMznd1Xe4oGv9J4mtztDpJleBm2ip3A8Z0ryw/7oGl+fV6SFNaUBXr
JkGcUgQC6pKf2ZEJLoHrsaQ4FoZoVcNK6/D6gkqeOQS9EXG9k4Tnsk1OgLlX0VX9
Q35Or+6FykHR0dv42CIPAPf/hkogulAopu/O29teSfUM5aDeUHmWpXkHs7MnqSUB
iWnc/p+7qFb8nFkYf5yZAWZnHDeJb36CrbrKZml47udE1RTtzH7r0HusxjanP/5L
+Dpf+MmVqc1FfUDiVst3ixkL1bCSBGAjpyTym+RvZaleIxpKR1o1j1QglVmoskg3
KMEFw3fE64TrLm8VSk1mXP2byJ6NwZDGLNw9JmuCtDpUO3riHOrG2GtqJxxscwf8
eZyQ7cLvEqJigvelXJlF+Tu/Y1xa9Nk6921Gm7wOzxhbkLHmR4IBVFUQ/j54v2lJ
OH7f+DQ1tkpEIL8BO5d0OGq/CU4le0v8XsgFzlxSLm3H0C8dNM9OXJV1CTxZm3DS
j591ZS05xjsgYJPUvfVCclPztpWtYzbcPP2DWGAdV5yUgnDyIsnsf1UMX3eDY8wb
UJ/f93gIqOOUcOxV3xfY15vFZ8YHV6SfPbUJwYFLt81xCmuPD0ogzTjzTOlCPIjz
VgKP3bygfCDyAe0lCnnx4ONsfMsc3N0/4FF1Q08KZDl6ieEa5JI8E3urSMlou1Aw
Q142tfTaoNsbn6eqn1YTPZ+XsEiQPIThxMRANKJTdRRKbzIkbCyqJNEczVDUXVDV
LsLwdqg+yJZPlW9RN298nrHuyX1kQtgwUyfX+Rp8ommOdQSQmTbq5hk+oWoU8Ueo
uEs0U/u9oudO4o5P7c9vXeAWXngD0e8jRpulbFHiG6LYFgyNK0RW3hqUEAtgh1Uv
x6ubCz3CdeqCQyRh0vI2R4LErzaqXGZBzviejB9WXGv22U2pWZebcBDSMSuPiUMh
gsRNIDdImhwcEwt1nLYLehygkEJKiTvALgo/f9AoD2sB5yx96a6yaqXy85k3w4ad
dDWv4/64GJO02Wu8+rS2nfCt0mnVz1JjwLQcflv9qbtR42Ud5ZQVayZ88FAMEVoI
5VtfUNN6qlljoFdTk0j9YCuS2DAQahk65fAcDqN6wtT5qruLDcQp5IeP6EsUS8ig
n28WD7dgs6GXbfstwVus2V3X81HGx1HwTctrzlIGnpMh1HMUoMWA8d6trnr2ohkq
ftXV5GrXmYxYfMOTp4Blheb0AKfz2g4y4ndkWuM3J+dBNpgeZ2WD19E3EOmSCjpu
hxgAdLmnUJHUFJHxc6P5Dlsnspeo0xDqAsOiqoTaVtSVzUfjBz7LVFgjfM7U22YP
spKnboyZiUB67sG/9w0lFaw3t+Uhqu9/Ve431RnNAKmmlAVfP/VKVL0T5fTDCXXf
shTaorgS4ZSBMO0PF/SCBg+tJA2Cm8uKGxBrP7MK6diMnV6iN9A1un0bMBDHjFiK
D/RTP1fIlPVblTXAi+E8bbwXR2gLDhICfgGPUgQJDOK8bGr6wh0L01rFA6vXb5kq
JbPgQNCRzT5PZPGxNAxERSqgxIDVvU1/CUdH2NE/DmfvPYR7wHH08U978U/nGNRp
DnN4f5WJl2WT46u3XNmiVIzG40NmzFxjcJ2i4Ux6n/hQykncNZ6CIwkjJOoMxcZX
N0U5TPY1tr8gjiLP0EoKBphu7cHWwnBtIGWc8ij6TZHwaboG7eh18rvTQ1TCDP6D
990hEMZ11Uig1MRnUDCw33OorJbvAcptAQ3AW03dnm69LkPq3FfQUnEpgrKt/otW
13zZYwcAtUrI3cF7kSvqf+jv4FlBH4duzdUOQUSBZnQ+666TsnGAGp1q/BHebxYK
rrOr2QY3nQEow4JpEy1tNatYZU9jFff7oTmo0jWX9VTVtXIt6MIy+vP2EzxLfai9
Bu1L0X3JWtZ26+1zjzpOez1sTil7jsJSiFc02Y/M8bTN9suxEcuv9+wbR7B5VB6B
iSb3ibybPorJn2XuI151vRs4KwJ91z0tNx59w3/l/vLcglL30AdM11Wm4WIUHaAc
VtiHxJ8ecXBb+kgZ6ZCFy2ouv9MafYPtobRoeQKQKu+i2G2AUbbi8fRVdM+2Tg0Z
pO4ZcOK3BEFlF+bVtOPONQqFnsoGrCQB+CzOsKiGgZ1cEBsHcKWaj1cFYtTnRnP7
eX/7n99BTJLstzpv94246IvpMlnFl4fXD8g9qW+m8gIn1o2iggOHbObJ1bM1VzXW
W3AzIRCuUF2wzT9JwRiWXu/cSmdZ5shyZiE6x7lZvq6KdUhA9i239WK7eYR+XdON
hvzkBT8c85DFKbB5zstLyUSXfG71oA3iNAUEPHJFBeIbNs7ZnsrmN9sTtQ5t+KKh
Xx3OD/G8YrcMPu+GB51dv9WXZEb8G371UsSsr3+L1YP1SCeQo0ciN6cJKNPLnD2i
LXuWXnqZuBKk0lp8Cnq6ssq5xbYIbQMgIMsSnd1txC5XAkoPI4XVSQjMahPBOoqz
c3i5BHQM4aGMU/Hb1D2VLjxmT7k8i3xPTni768BcOPtRXZBbJt7LzNWXY7LONhxc
oksgk8YxhbXEgn+kkbOmqxDUSbhA38FvMzE8UiV0Sh1cyZ9/KyoGFNiIkQrbCb1W
3bdLQaL49PLf2i0A9ANQBzvpXZ8aRqAUeoEgu+8YNoG/ElkewN16VIULbrRa4cgj
gIUPhNLOvjFCvcOTX6+KHw+gqPZz8/Lv5TG4VF2xvlUHmlUM3pqG5wXrC1a09sfq
fGA9qZx5GmHCIeUVKdk4UqdiZK6h6Lauxr7TrspWez8ErxO+IwVKnmXjnk9ly7sd
ROX8jiPgUpESBxi5l2GxbZSaFU544hGjL96iXQ0qb60Xf/8OJ/0bvGfcQUc8IBKp
etZgiU3wfVjnEVbnWgoVRCDRXKpir8n26MS7lKuEzXfg3E4xMh1NdClVr2CRhv6d
w1mEkSCFt1i5QJqxLA+HmZ8tOjjgbbHcAeH8mQEqBz6iGHHgIN/kUtEIRVIZdQaD
+ip4qybwqDZ0lrKVwfqnwPNfiJSonDcDaYLx0ZFdNEeJ2ByM6zXNIh6XD0h+wzeP
oMOGjWQQN8DQsRyQ6EBoDMlT0xnMk4NkJT2pjTMm83aJYRSsJUfoHH7hO8YxvpN/
sbkrYgeCqnqUDsxjfpDtQw4rVbudnfC0l3gDc04RbMG4jkQ9XzRODeJpqPgzwQel
Cs3I1vxyoBojxOLDzxJCL+R4+KaOXL3g6fzFQ72tp1u/r+C+Xv7XMBxfKivbA7Iv
2fXnj74e+7UAHGoT76MaI37icvXLj3PF1oQdZJWDXhYNZ7fug49p0GeYtdokqxE7
JxpJrutUSa71qMXKT87MxkqiM6oIP3CgdvnXvtTDGzGRVaFyw4KuLyP2kIckXgmA
0ss/CFq/TfDPsFJGCZTwAyADRmFYv4ycaTwwpdmB9gPjX8mjS74sMaruhDYSINiq
IP4VSmuxBiMIZPfiDWsF/RZhAwnqZ2sWlZly2HravwfZ3BGCuvxjg346594GUMZM
5cPQlnpZDVJ20usm/pWFV9N5iGT/5/q2cAchBx7AfuPWO0Dm7HrHHWNwT8y/H4ty
r9WuVUKDnczxj6cWT/u21Tf6QXB0WHDDajhqdhNz93S5HPObJxr1EZyU612qGRQa
R5ZUBEsl+3DfpoQTpQUtjFya7CTcACxHb6lEJGp8qAc206BOobhVEsExPwHECCFn
QieMKh4/xZeH4olhhfZfEzVyMN4PoQyL2xqgh9M3AP8vizuiLiG1pIFWUnPLSmtG
jFQjRLe8hJyVo0mTUXmz687+7T8YstGGa4UtViBHnkH9Fpm9AHit/kYkYSDOipGl
VD9WIFCH9GNdtWK986J6h6c5jX14A5pnET2g4xaI0EgTUoaQqheOLl68VMyifrSB
lGgd0W5dEMw0KtJpUmNzA1eH/mhNjQgxYdHy5t1f52YwgMC0SNRuzlHLBTrkvJ0G
oC/s+6uPKemkSUivw1rjvJNIr7Rm35pcB73aYZ4DECyJgOnV/D0hF3Xcri+Cm4/m
pdLWM8MVw5FG3Bdlq4s6+Y3polgbwun0mf/OlRPpL0NwNGdl9g0kOii04Ip191EM
RuU2fXgp06bzvD4S/T2bL4CprCmYhTojDXa1HGPDAAC6U1IlULDJAzc2n6SfG8rO
AnzxINgPxUpElvcz/uRveqzTZnB6CLwixUwDXg1FMkHb2EkMxoJoU+mMYlIXAJ4P
rZlJESqzW9QtHwzoiCuz2+XzQAcMT47HfH9WdrIoR6vFpuFC8fJxQA7X98wUzl5a
yP36rl8dx5QMgtr3pCJx/Uhu74IUWFP+lC7duwfkBlUaGmoMX//kuUegHTQgudiM
ZPUgIrRbnATzRsVVtgG7DrZQedjEOBs9MMqGz0TIAHzN+hYzbcFpheZC/R/63Y7e
RnJyaRxKJJ3pvzT0ZwQiNd6IkzlmMEPUBykem47Gbetu1822EwRvpFsRtm1zgbo7
NCjcXxEo5ZACDkvVtqrFpkirEVBxfs9dKbEh3oQYpjAI4YU+PriKQ0JN/MA4fcMm
/VNhkc0v1ujPopyAh+pNQVu6x7aT0raa+yfqPyVbLsmXDD6zKQXm+fcmNDcUNj4P
+xg734joIGYL8ibJR2/6JC4Qohmnp7iWVnA8cz/a1AThFiQk6E/pCz+WoO8bLfVW
4/wGvRTmT1hMPBq06gTC182jvjSPOAmr74CFu7Q+5de3/7RkOw90F/4sF4kv+F/e
K25SvIwExurCxZI6+KPWO6vk8itY+Myj4FYJ4tB9PTmAvaiTIYdHbIYXaf0w8QAd
Nnko9JqeA7kD0pMckjqhAsAaEKcd5bC4HDHRBt7aq5wreLzJs5H0Xqonxz8B3YrC
F9y+iULHggPf+tTl3lNlL0ibil+Iycwo+NH3qcGEKKmYu7wzk3Z3hUcWJrp9+zM2
UE3+fuW0yaVAfmJ6d7qI8WMT3fjuA2vs069/+2nbrCZs7MQ4pp8W9ibExgnAAxat
JvHb/ZbxuUk+F2t9wqBSgdux1P4HGlXKPPCgdeVtYK90owkMih8SaPwzI4woSefD
Y9PMyF3HfER91ZkuipartuiBeTynH+oxmhmnj/3sBtG8/7ROsjZlfLoYXCnFihvF
dNdH8jptaXJe29yUeyeZjPJmSOV9bDFZHUPcLYWp6cQyqAGUKDNYMbRCTO1YWfJd
2ildQKGu3+b32PAhTwNXgJMiCk8w4ETg/hjK+1i+muSvzdEO2+gBvLnGpozvbTNT
SI//mZKrSJ+an7mxnViC9ROmtM+tIhHqlrF1mf+iWC7ohW0TItJ42mQW9MegYQ6/
mRHJuJlLQFbDCsBGMKtLYGepVjoiM7SBxWhdER13XnuX5OoAtAxO7EMj0s1K0Vxf
SsB6uHGZgxU0nt/Xib4OxL9kbUi5fty7yOxuf5taNnTSWwtproAKYdtApy1HVwTR
/ce8P/q71jqfb09c9CA+/jAmsBtj4tWIqsAztjvmpZ5VqSh3w9F/Kzs8/k+f3ByG
g/4sVDumuGT6LNYXGnQnkuMkLwDvYZN3Wtnn9XqPwy8MJPwpPRSwzprx/IohuCss
uSyir5ljlk2AQmDxLoTEi5UQdwGjLSCngbEsrJj2Xmco4fQqh0upwgW8FwgKpZIq
poXEDvEBPpq7Th1NEwfwTPdXYCpBiqh0dNUdadRcEmGxKHEyTZ/18FqZT0Y0ow+K
vDKmTMunnGxd9AqWVETLXurIjG8adqpjOP8kmomd2gFAQj+DabHlLv5hIJyw37KJ
fBMA0JdW2q3EZHjIAHonF5xzli6NZhVpoyzMqty54Co++tXWCt9AQ6nRxfUiu15y
AYBEcAW9NBEsp2meU/H/QAfFWqJ1NkCPcoJYSa8pClAJ2vYHMzQIp1HB+Si3cAtg
gchor0D3HBi7X+1c9cKjAxD0UrNflj9kaTTz3fpcPc3m4E4VLJodyn6P32pqZsy6
RypkpW1SlnCnui35v/LFcTb/nBI/OxlLYISCNAq2zWarxzMLtlE2C6V3Evy4QnVn
6g/UOVq1ptAaJFvOXIpLx8KmbM+Hkz+oRudGHnU+XuFd8e0xTo+4ZawbU2vHOC+e
/H73g6pi1H62CUj6430Yg9i+iKRzsw7Sa8d7621FQb15eyJ2I132vIbPTMIX6Bph
+KbEZaR0BzXC+2qguiq4qd1KKEBmE20l6OqXmEsibDVkWjBoQWOiWf8YlYJtdJQY
MXnFxp4Q3By5kBmGk6zbNLm3DPL4yccpMzF+RboJvbSgLbuAkZAJk97QmXD+Iogy
POM+PYHGaC2ZHz61zPZGapGuT+9Ig9eEsx7p0XXONwyRcPspIPYrhMEWpQfJ+RlJ
Oji70zAi4dVVZWwmU4EZKJLT/RETEb1lK1gzMprZZDjzCJBpgLZcfBi6o9xanQgH
Kdxja1aWAa2S7meJhjRQOXpZQaXWKzYHonVr7UlvzsKwqvTAgyLLuVDfhW5T804X
oeorllwrgDsb5JVILHnUWjuksD8hYFM392qFuU75TsFbkQCpYdaPnGaujAfgLVS1
f5mdsdWwGwg/vBgGppZxVYtsirgw5IOjRRPGWQpoSwcHyXAZB9virNgZaCsXtaHD
B8c41IpoDiBS1FKok2bCcM5kLb7OmgaV5OEF6ANWD7BO/8sttl7BCTNoGszUJPtw
mAQCOM0pcp0jbSvFuLRCx8k9GRXkTXffYid3k28tdMffpRZEkNIZ5yVoQ0onkKTR
Sr+tS/3ExBe4p6sSrnEpEsE/q1m81ygvJc7RrkNuQHc27kJMlFVxlxLirjOMSFpq
q4Y3gQ6DEF4PwxFEj7qnGiF1w9mNyqGmoEK9LCoH+TQ94L3AXGH+I7CgEv70TeYh
k9oFXVR+tmAIiubFXK17IXUwZsU8lVmqFP8VgSWfsOIcE8QnPawdGV589r1OB0+a
t+zxCiH4VuKsLaX7OSieiA7k8V+1uZKJOf5/op/+5Tl6DrMzEgaZB9LJNMGasfYP
kvpTbgJF0RM2JRsvTfX4mI4/jQNFlz3ZP6SiEh2wn2IRn/u0xczbOrgVksXgWfSI
mqAt+F7mddoNseF/89fc/6jTnsvW6sTYU0crioy5TMCVDgy6mkrIzEYnQNTRcK8S
AglmT5BVbBCIWpjvmrfIc5M0x++vFEGDUrklf8GtRJJPq1TYNYpQdzDguVf+GWyb
K6yhebXcFxQsFJoff1cPJzGQwYvgwYT8JfPbypbLyynTugbSgtdxNSqKxQPZl9ek
XUd9HkJMo9qzhx0+SvqXo1hcuykHhxuFwvwVDhR6uHAByRxpUcJ6jXPwv1G4+GnC
0txkkSYn6SeyqfE2sMVpW3ygq2P40C0mF5ccBOY2dzMoCiX58SW9mfKkgDsnuVdc
zSiCmY9gXTc5UiCxrOUtvKH1y68X742AlCf0SfTr3Abgm/7KPJXTuL7spNsqinCs
Yq1yIdgPo0mL7fm15qDXaxlI3OtgdvPOeJglU9IhYBLYmbWJNaAUmMIHq6PR8k1h
QEMgOzurO/NNzNlQe8dHvJm6GXvQ08TgXZsj+2vpbM7qTyeu7QbOwVMtQ+Uux6qY
jniQwYcDF3pBjDonmEHy6OYE9KDdsRJo/RWHOg0NBOZGimEX7TcKZgsDfgCWgh4r
P2Yq2Vo0QX0YWs9h/DfhFedBm2t+mCvNTHrekrBVTkURIqipE1FXOiRWgFF0p1g+
RwwdYxh0A7lPUDAJNxvEoFqbgHtGUFCap7q1DZbmZgrCdKaHNW3ud5H1X75iawP0
09QsNi/J1jMaFQoEPQX7seZC6xdctOIKJHTk/3rXc3XUwuulD5CKA36G0/I0d5By
bG8UZVLmlUFaHDGwzE8Ah1HUY6MMI9SoRAyCiSMJtdWqKf+QrIYZ6t4M0WxsEuq1
5BoZKCDXZM/BowWSHR6SKTYFlxfTEzBTNcE0bgn8Zk7Kpwzv9I0Xp505G/yKIC2x
dyWsyFd3E0tyZMpvyoiKnUF9wlvIzuUy4BL7St9QPJltuFn0CeRKui91cBUl3UNf
FcMdYPntlU0vrmwAqc9IEeZ8xPkuT+XtgX896mHzWtKOrpcxFlTXjT4isP3fO4Au
tFxd8c9AGN0X8KQVSjSokkLLSJSOzF/npBfQEOfq589qsS4ptgEJ6t6dj+c7pUKl
QjYhxR75dmk5RRvCuGA/lAWXPdqx0iW3RyocVfn0g/+Zcy6YAAJxfLSZd0Fp6p9s
8VIGbzDxNgiPA8/QAUV9sBENh7Mpv3IWBVUttLJBKJgyAnlNqqfjKmNIpCpraXWF
zfKu5cihX0WfXQ1PwaODkNeSkjLWAwypF+HhZDGuqHp+TMqfMGMdTYSiEq+Y1Xdr
l5ZxS2oK5BqX8m0lnXLfqWGXDfdY/qLPaUnS83q5CEJXuTVEdjCiZQuXZnjbXrIK
EtJozhnmg2ImBeVO/CNEp04qOWDXC4I4bSqhPIGAgXnogz1eMNS5xH5mDfVhv6Qk
QLt1ZzTb6VYZ3tpLL6w37IDKHRuMiULSJMrpWo15d5QzMYje3NSpRWvJGDE5P220
KRss/mNNfUPzXBJdRVu6b0XQbEu6KBWZt+2CuOZ4xZb/yDFlVawjO3wMVGCGynoS
Lw5IEjNZuIvWKCqRphqpt+28stjNyiMHW8k1X2w9PdzbXbQulLg5rK0sBvkC2/Vw
xB+WyE9vg2MrCusYdXo8oTOlQ7OYENfcIaib33JVItY4K30f94zE7j58RhNw7vvY
jek5schdoJsEF58Fh5HoCGbGcKTSiZ8L+k0jgRcfOvHMhCmiE9gHDQoAc3nU6IU9
Ac4lrhTVKKF1Xwfk5vd8a38iyNKAHz7w0YCrahoyA7aMfVBKUG1X3DhDVYiF9CiB
niWoDDyiUSV8WZyCBFuOW49TpJyJs1sVr56xbJQX/FzJJIduHPZC35fcohkZkPOm
IpdG3BC/3QKGbCnEX13JZzKi+jIbctRx0yvtSnkgycy7apcW+u8i8wcPi2UnKlqK
S8gzfXigskQOWKTM1/HRkRggMa8zzmoBFhcgifS5kYfCx79rCpLKJoH6w6fcsOMc
BsEDcziu9owTbyjjeNguk5AfjSdGYuWm/0HapgWkHTgmavfeTk2Z9gWRonxmY2iB
aPaTntKKLPATrF2IVHpHdwH9PdGarmzqT9s1J2A4bpLGLhgXTN2kMZ5+yvhOOiSx
ojOiA8xLMlCvoUuZueV13GZQWafzuDFbU+/QKl5CUxebZdyHSZ/ms8+TeWa8/pb2
PSPtLuJmzFHlFAqRO90ijO8biBNhrC4LUfyatqi04zWMm9X3VgZxz9O/WXzF5Vwl
W0fsU6SGcXdyNSB0orXQ7feWzw/zOXpcxf5I6MGcfttHKg/d1Y587bzgvQ0yeBVJ
W1riQHrsfbih6gXRA2uaOp241fimc+2tnwWphiyVJP9T+QY8bqoUBRqDYs4nu162
wHkdpz2HkKST/yBRUADGx9BK0y2ntfJMUbJXYjoAKxhRpAktyycM4TX7a0foHvHM
UMWZ2IaqoczRpiZU4dToU/8q2NyW6X5rBTVc7MxUJMrbe53mMbkNX3+xVSOB34aR
nrGGBGr2NkGFO/P+8kHUDSSjkAyXtMUDzut07XX9nYNMEkUySQ0lSHZZXciF2X5t
1avT6Hjrrjs74rwBG0muhghUI9onltLPLqDZFQje/TIiM/4Pvikp7eheMQdVyDvq
qbJqdKn5fqdq3+o7cdX+KJJNjCoHvjlIWqoYlVuMBDF5oB3/3XDjU4k/HfGdUOPg
atJ6RoBdaigIIY5VphMKZ3hzWpitGdQG/JygVeq1Lx5UKtyGDfUjIilQignjrw8m
frl63y7qVLQkI5T+CIBSjGAvhPBJDVrN7Eev0hMhUSBk334p10Cg8GTGRKaR4MbS
B17xkFaqFNMVpGPHi1rtdWQ3EUk0hRXWpaLDL5IUIklKZHfYJUC4LOqTWgbbmrlu
wZbeBHC0T0CvckUA6EExHYjnTJ3DEuEo8YEfCGrrqwsNoGnVNLCYcRWRgCXQskpW
GHeCETQMwfabrBGSp0VftctUEtN9SJjHizkgqdoem0NAfXt+NK0mp06gCT8odwDX
bfXxM6Mxtu0pjV7u3l43v/h+zTcvqtvS/65okWGQUGE6Uebpyx+X2M1wLkPI8qy0
BWhQNLG5irvrEV0dQopcXG1Fj+1mCGj0Hdm2UbvQYh7lzVoS5cH+XJSAzvudbPXJ
iBYI1shnE1fWixjLbxui4pDIMljD88S9I4Qy8ivLRLLdrerHoMj+Zac4V0g/Qeaz
Za3pLBoRa4QL2rhLR8ihoZg++o3ImqS099IYyec0U2ZF1dXaTPysaaVXKIelsmNP
f994xq1jAKFpYyemGLPlukl924M8dfXMPWf5Jk1glB+gBmJ4oXR4k5wqQFzSQpKv
AP9vv58hiBWHwm9Ls+VdziBJ/eHzyMGOKV1m43ht9J9oXPSyVeEVMXQ6wxEgEmXB
Ops6FjIPSzwv9uuTrguWAVCJ4LMVObjYN7b4pPvHpc5kzHE5iNsM70RZ3HlTe+tX
CI2JI/ej/rAlA+dFFm8CcXsoqKolrYs4zpo1yUuVnGvFTnKa9kiJ1IcDv6jWogh+
o7nGWht//5YLi5h7U9PoNcNao+DztRBxtrUKi7hZGnyr0/0fvEwjGGUITFwZ6Dvn
XhMKUkrwNm/7xK2vYsPqz76ceK1hDRF24AKNidiLU1Yq6iy4M8XrSpgyfAzrR8bA
ll5FrEfCdS9wkgJICSQhop9p7bCqMLY+6t3eo/Kh2IuOYWRfyFrPwZpj6t/9epcD
rdVrMLFbnd7GxXldRYtUSTb2aHaL9QESOtoyGaCSDa7wX5psZHfx3KJuWeM2AOqm
WCkSLIcylhONfbCkcEUo7s4R/WMGv8hHPWpsmR/HmKZEsrkXNVux2qZBENm/47Hh
Dc+1u5RPySGxsog0PzPPTZWMTgfL8ZxxXDTWpycBSvL9RI1xYNnAw8UbbhdNKz+t
GF3KuPBqwnPE+z0HUlU2B6SZOEBrDFNrB5oMP31AE1TFNtqy65mY2xgLqrZAeJWS
7F+1/5YBUn/VzS0LmChvOnwQlaK+fUBC3CXiBv/NN25DvnT07dL0UxLY3HOvJiJO
QsDAC4uyzCUQRCbCu85zvsik4uB0pD12PJjNMr5jugxZ2+Sd6b4AJmNkvJggUaxW
2hVzKQOzSvtCX7TiMVpOf+VRagyn+dPGqgXOHfPju98oQ30IynD+tMcA7/DsSEXk
CARej0mkWJM6og1qfS1dJl+GOJS5x9yy4QQTndyLQaNWQeh/NgPY+gF0jMo/4ALM
wnDtXXCZ3V1joIJREvmHvQplJEebm93IZrDpJ26cgggXXutB9CGjtcpnWdfsQEMr
3+WvZi8JQRn5qhVBCk1PuHh4Bf6jIwM7+0fjolQXqdW3+nsQAC+OpiLMuZ0P/zRl
vwLHl4Xk0EJpAdJERtu2Mj3s3TpPMlI7ntYNRqatpnSMM507d9y8bzc9WhkCoPpb
Z2MhxDH2Jje2LIwqzI3VN7pV2L3OVU55LhZmUWD0mVb/Xs6/5re9xdTxuE8hScSj
y84mcBoyCd00CPMTDBJhFJYs6PB0YozN+sGTRp+CXsB73LO5Cqk4A3UMHhN79s1h
9+EJ7SjxT8OpdeWXmTtHKZATrtpJZ30kIWnnbeGHjWjN+S9drmgiVmMas3auYDc9
MKn65ec+rPqB8PPNcs3GU+46U+Bu1q8qY8JFHYxCAKbKW16uot0AUD262W7UT54H
fM3sFykOchpCEPyfxKW8nGiygEZJM2U5yVpb8Ma6IZiW9GRF5osD8wmwgFPCxoUR
KxL+h9f8yuW0aIoTarBtAnQ8A8dCK85A459iz1lcw/Gj0d152tfgYlnXTYo4y3v6
1R98hSuyDj+/N1UGMwTcfsZai4asBo19PnPQgImAguFY4NakDYenDONx6bSXC/fP
r+XNA9Rr9TpcQKG86lZObS+5PLfyk87IJ84HtlhactwDDboWvI2iIyQwZ7ahyFJv
aJ1gP6EJOd5ixJnB+QgoTGFM9NY2u4b4AgJRXzSdLc8hBWj3dJxNYkSaqs+l3Bcf
J0lFSaUINnqtRaPTe+g+sD2D32XxzTHbdzTm+fBbC0Z6WQRaxQZMJQEXOMsPb7Wd
ANIV0ICupUg2cp22RIbm4m4J4BeW5a3Zu+rW7AoRbTStFo+0Y7PiQMMnpe8Y+pBi
0Jd9Oa81CtkAblddO2DAGmsoIWLwSNKo6p7HP5nIGRxERI9OJ54SKNh9FeRKEGMJ
yVUJMUtCh0dca4Xo65YHagOd+GFz4OctR/Lhnevo7/sLY0ACpXtS4YdPVKFJjXcP
+gKYHNw7FpIyierhP4OAFPpCqZItYwqqvfpCjnL1SRRlkJ8lEH0V/QnTXgnpyQFM
iDvDFIGLmilGstzZNcotQoubbqZdaWwpUmzOgvpwwX45FAfTxEguyL3DJqYijpKn
hL1e1vcip0Qy8Q9iuzYluHS3M9oegwxdbicnu+1XUEm/FshOYgDSCGjMjwiSrfFo
Ot1b2tcE51MbhZvT/AQi3ZSianThz18YD1iG2RTmJXJcia64ehqfBZQ/v5DJYXoR
NfbqDirkdjsgKswq4/PPahkoPwcqAud2CmS1l+0C6LD+RtaUE8Hm34Zdztm1pBUA
wqmDlvNgZYoA4BCyGbhPGrPBJW85RQZ35itk9GjOyL7MYzR8ZBR3PE1v7oPRa21e
97Qwoy/UA7zNiD38tyAPba9jZD1pkotg/8V4+VU2+7bkEY1CnhR4f398e7SAZ1OO
+PqSPQrRcMUb69WGsZRAo43RFkc2MzcMcFVxogrF29VdtU8sW6RisU3l82FGT4Gw
ux2tA2HcvcchohRd2QFuXJSRIyO3t3BGztlaIYxlRnhNO+p4q+hwMTqO9lgfYLvl
1RcbmsX4RBvncAwHElCxZM9nG3XucjxH43T5cYqiQq0/F/ZhK78JwSRsDef+JCyu
lo08q7saVNu7GuAXC15vObIOK4MLWdf5PXoIjbjbB5V3TX/RzD2QdS+bb+HcjxDP
u6T9goRipozgMCFJlIFIKux4oAOIMX7id1XRJ48svR5C/upsZexVkQzN3ZPrmlqL
4HXf3ZxP2EIQRbbjgJ061j+hsV5UgMSCL7VSIndGnM0GXqu42B2gFo6p0djgCcEm
PmUdi2tKlFC01A7Xu1cd0BPn6MKjGI/wTswlqnwmA++r7JKTVIG0BqqR4YxXAqfC
L/I5qZ702af9d/evXBNjMfs9dz0kvCRLd6xemujw3RQEAqd82554gIwJfmg1g8OR
X3tePWqOtbD2iZAocCxOfapqbMz8m1dpaDZT1vHOrTVaYfnWUHMNGhUR0XD7HtXG
6pFt2d4CbZf1YQIo03219HqMf8MoupejbHBeaxP1AbTYMndl2YWlREsmke0Hj2Ih
HDBItVybYGXr1y+VRwNWOT0tfQjUB2BLcuJpleNFGKizvEV/danaXw5sVoYt5WJG
mPiwSk+44J5yHU3EwCvj8tOaMZPuphSDnJWi4rWN3AaktUVCxu0f5U0FHcXgRBmQ
9fHlX34bSmRyqp1+tu3YOwmK6wEwK8OkeHhwJigF6oOz9IokY1Jr0FQx1PTQpT8B
Rj0w4jwTNTrpHAHmBMO2ZQ3pYEVbJZvqr6UDBHFrGJgswFQGGn30xojKMhB5TGSJ
t15LqoEBgbdqRPqjfomtAJJRdLym2WZCd2PvzBo/yD4Hh7obFznLPFPJDNcmafeQ
1+HfEwR1zJgciltRlnoR1lyGLNSjA8OBtyMaMI1rfFY9wWK3ZsNuWZw2ZygG0qUO
FENXH5U3SJu3dny0AV2DP/6klGyR4vAyU5fMC0CDRedFpHmQtwoGMrJwoZYS/egk
Mtaurw8AelOky+1Vc5vj4ewU7ITSIc5eZy/yxXi1g57qdV4kye1ham2nShMqy6UD
vghTn8614ictDF3e9WstwYF27oV2eItGPjtEbYaywGUoWkfE+f9qNg2gjpbk8+Q6
WpQlxxWFegR4cr7gOySLUjYtw7rlc/eJXQ6IuIW1n3E3nPFMMI9jlbNY01WxhrDJ
jaJILLgW5YveLhgZnqYtlpJezHhvr+FWkynWDW7PMRGNARAclbU80uoBih4RoHMM
EASUeVGSmwh4RflK6PUD1NX+nBT9LeLkT4zOwOJ9N/CDd/FP9vjDg4VaM+J2lJK5
WoqCKRZdCyVzUubiwX3HaVvisvNXN42pt7omFUDSbCeDohvY+zJxC1Bi3vppuRVC
ZbCJlvGm8rHZGieAS5CfB07P/zcOvCFnmGr7fjdnkrKemr2RD6IVU8Urn6U/HE2c
EWHm4esgnKJ28Aso2SnxGNP/AVCtcvuhx/egbL6grZGilv7lHkYnF024gX5Ctu7N
2h1ZbYb+vmKo40MnLwWB36HpC7rh4jeeGWrKbdp88KBNEjBsskcXk2g3ZwUNVqPc
49nB6bDhrK9wfv6d+AFD7scKsjN2dv+FsfsSEXq8HD/BuMGiIj+9oUhltBkskbTS
thcg6f4Zi1iHUnw+8VK9PmKAKxfFclUJkW+dc6OV9KNJceP4Cw82wzopP42xbio2
XIg6h1X/fQRT4ZdfN5X/D7ZrRdIfVM3Z/2hGH3ZCHJOVEgyRoAS0Ci4zbzPTR6VB
FBJ3SSnwtGDhr2PDggT2JLaHifJsOON8e+5z4KS0Osj60engxzLwRl9IEgQEdVYI
8bphDyWDdagQ4BD/MMMXyc9FN6wPKKadh+A8Dwemd9K6WkrJ0Jy2d69tGfHtQEwX
NU7Yxrg+06qMd1H+JxUz9dmm8mS07N57dpgYihxICVQepbncIGTHdvpeVETShs1I
R+cJ7nbyrWsEU7NMtP0RJZ0ZGVr7poTdcgxMsoDxNem0jRgyLt351t8X0eII1MTT
iVWpsAl0VgfPzy7diNLfKDC8N0K9QojqIHXL0UUha2BF8EB5orN4KppIOAo/51XY
CAkfAJz0T+uUtTFu13A2LuNlPgV6poFVta2L0lrDIr2DDr59bRoOxNkXWAAM7/Wm
9AymimzXQNnSLatJwhB+GqYjRAk1JZUqGH+poRgYSpWPrdgeXET47TEQPhcBoOXW
36IO0Xf6oqbYgrd0bRSKJm8o4c+6CL1/cIvcJH7m2cBx3AJQshl8eQuWjlDr/tww
sWdf7cTHNIGAFsSmluPQVpjGErUOcFzxn8M14oNLrW9dk5betaKdYq8eb0on2ycr
LO2/pLmy+hJdII5WElHtmQ6HrxH7r3+SzR8++ILmH/O+Dex92Cj0DUdnegpMXWZH
wcOvNPAg6L3WkDWVIcCr9EFSZ65xCN2R7vYwUGLct/B0wiV7Q0JA1L8HBfH5/vSF
kInJ4vJO6pceBq04epcgEL+21k9lvMmpjkbzCQJBNXBkVWxeMoYuAWt0exf2aT1k
uFUI1XwMgzps9lnl/aVYG+yiD7HKlgIZ1ZDoJ4yOcUiWnk/Mv2LOOOLFqYFfWAH3
kpd5ynWM/nUVPHoIXnup1J53JWMRwDpf1o7y1RMqmwdpgy8cDoYOU9Z3vVFWAMTX
Vh/mWhebhWeKjVYHIjX7FibhnN1lnl8hQPMZAQtXXKSxT1yvb4qPTe91ZpQgZgKu
RKORPRsZXm/nHO1gdsuYTB31njV6ySpuZWCxkkcRvuSmiojUnnFOoufI1QB6LgPg
lJwDqjPmRXGNcsiOapJ7M7t2TdVVTTCwAqNqewH3qkVujjViF4lDBjn4IB/XoKBj
iAf4Fhi4gxamXt0chMDQDuSfkJ7DK7kQPRtPwL6p8PlWYPtEQvWnR94pJRYl6xmF
06WdXRDtjduX8k9YYBZ6x41fA1FN1gt0wD+8ctPWJ19RIoiFxa01c6Taq/INd4a1
TZYUAFb9MUPfuZ/7vCVDhmRLiOOkMprXLXdvQEgu0mutmsBnSf4RkSR7fsmZLA4w
fPtseG3ZnB8WfJr3XUQAU1nQv2l245fJvRhAfgRLsUGmZkBASNGGpX1XMzBgBv8Z
82ntpKnDssqyUzVJGNmrZ1gdzZukXJ7SysNXbEPfkg340SJvf32vvILxK4goasEa
xxJRo5DAZ/zEkNi3dD3d0ezgbaY9HPHDHtTWkWrF0/bbrcEWfB9Yzzi9XwPR4mNq
0h7mm6iJJb6HrTgd5MN3QjyWlMieQfORzegnRaAM8Nplok/5Ht/etEOZQ5sARmV8
TrIQUBXgSNUgHwRlA+QWer1S/unvVa53U7hlQORFgpC8f0F5HneBlF7l7jBR9TQq
AQJ8t8Sg9p62ytbSFzDsP/eFRktO1BAxqzMYpFtttOZSHZMmaNDME9vMvAYdapXo
qxc+yDkGqhPI9lT1yWl9zqdUsTrVmYKhNc1Kgm4JhAN+naQ36dA7VSjNpa/3+kaS
k9tl0eijnPQSf2eRxlM7kOYeg10i7UKfBlSy4Msu7KrdORuReoZad4Kkrwlpzgqf
fzwYteXnbrbiNYcUyhqaHkgKf7Jb6BN29jwHG96pY7b68a5fBoKztoWJUW/EaC5z
TWTxCyQ1fw7cba/L8t8v6IbAmIIo+bMFOhRiCQkvsVoSXPcrPJTDi+K2/pIZOml1
5i4x6Zl/ZyC/Ee403SUkQXETaNMYKow4pT6iCmMKiThAi6WqcEfhMcmxiKaki/yz
ZoBIqFicObG0LNaWhmw4V0UC62onJfi112NVtxUIruE4q+2BouQ5tRGSyP94J2MK
ElKN5oTazKbgvcngDnYynGbCJJN67q8ffE9bJu2v63LfS/zWiECtIVSLgt8Roypy
YNm76RHonN78r7i9KVFITC228EqkMKHP8nnQEtD6LQxUZx/ORE8pWhXTyOuaPkNJ
RutfjxC64y/W43Mo6rMmHBF6oXxOYfKwwuQmvEoTIlhI3QCdA3ji9uh8z+13ThjK
Ep/9XUDq1EeNO923IRfzVrtll0SsZu0GPQyvJATOQ1Q/MDgwTKfOHJhKPGfbdB6a
M2vQRBGs5p1QbxmxExCufyZnH1Cp2mheHA4o+SjVUWZ9j3LkbkCnOtV3vEiBpuUn
uNuBRoiG243YdHI//Q8/c5FjWL0zanR4rEm8bhDhtg9JkIaY1ktIP/NQsKO/TzQL
sDUKFtvnB4iWOjCcgohPe3lwFQ1y8Eea+pVWC88ZjIKjG7Sim8srx6RrgZYPdTfT
57V0QBgRNi68ey5bmg52pqEQlerHBukTGooWODAbCPFfeWb/6esKYT+qOC0ifMpX
eeULGsyNqX9MxdRhmxSaQdwTRHFlATxCyD6eVEOzRCeCoypDX7DzrzCH1YJbXofh
w0VQCxdUXQfttZszv8YRZhDtdeSk/ueUpbNUTuZ5ip2goV12zIgvQ+wB72ENEFs7
jfzE1JrxpVJkwvjLjEhaAWbOWHXXn9HaFYZv+RhcvJJR+35u8rZJ3osWH+BDFOwG
ODHQafEM+QLFr+pbb5o6a0mZArgYuLUza8QRdwujpq2MGxAOJ0MsAxeESSyfOink
/JVaN5EAYsHkTpZliEvqhf8Qu7FzMRix27kb/8/lDA4G/Cl7h+CczVSz73uqs6A1
J217dR68ouZNB+sMEZ9xdwYQ/grhF6xn/YEHjjyKwM7J1tnkSN40VtZzVQrAFJnr
cj9jEgE2LtDpdlmRSk4ZeTsseKRray9IP87seIuOnmk4e6egHDAQz99IUr4gjpph
LikbnWAAfwnpK6i1wBjL2+XfTBR8i4rQsalbfATnkPKw26JF4SkjRuIR6842SHNv
+vJSGCnr2Hwq5Sow8uC6J6hiJzHf7mA9G6+zsd7EdNf+xMLzrf/vw71DaglrqXm7
uGDuySkOubpJkQfLWcmiQNv3MiWfKHTjpa1vxaa+tzSfJ9BqKNd8eYmwaJUNZzbt
L59xs/dadP5qxghVPFZtI64CqQi5mCXfB9LYjDllhhYvlWlyXM6RPMYjRXRw7MyT
Jp/As9OluyZfaYedrMhHftRIbDQS7vl+37dQTyEmDVrp8GCRHtCTEUmsfwzA+WfB
QNkL6sSj8YKvKRCUj8soJ8X+N+NFQFtLhmEpIo60LtYaJB2Yb+n4fAZ94M7c4GSd
PF2mPdVSCDuMbfaQ/tEMLxPkFsQVwJAjWw4UHYAJ01FCxfW3xrxqBNI6CFaTvtLG
T66NREu1/9y6DEtU5bJOuNKusypA2ybl/leePxq9pDdt1Jq4VbBtu04OQdeL41D7
q9KGx9ssBldWoqckqHow/5H/2CvF92PnQtaR6EZFGaeH5X+PeMDHLtuSQwTHDq4p
BEs5pFjRlGwMoyAvhZy5DcFIgrWxXfVNy1ualKUfhls/4b4ikHHyIAYiGQCulLKe
S4eiGkdhPV+FRxQ1iblDvr2BsiVJ1+r0Ku8rUFGRtYtQL81jK8gtIL1aa6VoOwFd
OHg/ukGLZi4qsvqzu+U3Ps+QQgUFVRuYTWBsKbUfzSxLAagKNZfLHlhRpPWdEFQS
uhDNl+Z/xN+Z74V0mD5ZEg5JfV282zMvbyy8qvgnd+ccdv6zGP2JUKtSlYMu1wnm
RbSEd7K+7bV3u/m0dubM7e3UasB8xyiDSbG8FOoa8BGXsOfHxfFEMnwmGQXEJcLC
ZHKh9YpLV17/21VsQePoC7VblmTXyMVDXdL8E4TahErOWMpx1c6Eo2YiK1MC+v1o
g5OYF3H1z5ZjacRfSl/b5vVuStix9vfr5b5bbqm7d+bb5DaY+aWxqscI9DQsQ4nC
pyCq3qnS0EjgrG4gmLb3bkhcxuDkMfK+w9ryPlYxMaPA0HJ1eQjvf3cL7evV4XBf
QpPCsOZ2HigELEsOnSnDpSqzzOsKOc0ZFMTQgFPq7+rcgxV6sjzEvLcmVrvti8aM
TXcG5B+CtVxVLLhVmfWrnIQKAG6dMy9sunYnfAGlPTK+YTk93c1Y8loZD8RpSllH
+VzPcVdwnuRjFVn26luOgHkWFC3IWNPVnun8kkq2kM2J9qMWLhWYja2zgxyhmEen
Yul3BMVaPwWjoK9NPXfgZ0QJQcOrDaalfVo2sKqGSZgtjgk2pU5KVW7wS3wwKhCA
mHM3z3mZqRZCmOHxf/SGWaEBtN23xQxwO2o+nNy1NFFRIvZADxWCPJXri98iIcgm
XSyn4Utd6VqEULDUVXF5TP7a9W9EuY8Kjh3QfBfyxrUvhNmmgvSQiCKlrF0nL9EQ
WmqVx/8lN2IXmFk3XvtlBmBDsb5rYAZddv92ZsDXJOwaKsTQRw8HTZJplXBE36Mh
vmNAMHimxbhD6wOVYg1wxcRMAr0mi0pBKbKs2U9VrEbM9mbzUZCGdI3B+oxeDsOx
ZSO/ihoXOTlGkIbZFTy1EMZd31//ZfRuZo+bSTFXz6mhuxDe9DjF6M0uFT3LAjC2
ZJj8q9NGEZVNGa1bXs8R90IyZemscbRzoYDcO0jgzeseqHgqSDfi1iCHpMYrBbFY
4rNL38e105NoY7mZyiJqvTwm2W977/givr3JTDU6UY72kcJRsaOU5Oh3bR7isAYq
jMFazwIVJfINRGqaBTXDWborHnnwUB2lLZGadeYqm6rgWANBIu/BnCyjMAaNLLfy
dsF+SdGxJ1yfFE5vxMkE+3iMjf0y28+K+wILjwVktNuP7xAhGE8TsBYz/Lf9J14e
dlj4JkKfD/RqG5zQ9nocjL3bhx1iAgRbBnht2Eamik5NrQlaFGFfkFepM4MvM/K5
ch8LrlFmCWvKuwmQHRQBGrSPfrgyrTi5Mihv+mRuCEtlBL/edlzlKyNsySpe9wBl
EAvutunx3yK1JQ9Z04/2sYbxWDMOzevd1WiHMVA9EN/mboNTc2BrVfY5ZX5PF3qu
zP0qpi1O1LMJj3qwfybvMSEyvn/448lDtoRnV2HsOHKX0KUB8L9P7KTIrWJZNRoB
4otEmLFfR7awFR7fvfFvmfMDNw9ymmdWAQH3QgOH3vB+VYWaf7SwKCTgrXT7509D
pEjtt0FA91PjRCUHHw8BsbaZqLscg2Ps1MxpyWIYLG74AleEQDdXCDCKDnlOnPhc
ZOT/9UPhzN9xDMciN4cr8dax2/2VR0xaKlx0Qua8ZKbQnR7vpBxoIRMUUlMKbHKS
V7xo/AOIXLEsmRSy7UdOAeTVKkhB1Xe47GSkhgpdu1itdpk7WUzgAszNhGbU3jZP
fNv0DcRVILYiyh4lbzSICeD0yqrnYT2zX44F5R1wiiZq/9GwT8ldgSkxPEC7zL+O
zjAuJvLEzGLbZz+YdmK+LWOn0M7NsfEjHnuN9XCvVZ0PVUXV1Ko9UKL+TqozeI7z
J+BAwdClfUB6gchRtHYNxpssoS9LRzGPbH0x//V56zZ7Zt7snwpOFkHCKThMvLMF
LZ4EjJ7xXgMOdmUVEXJQkoN4+FW27EYJbU9RNAhYZ6RUMWQ+ke56+rgxUMeq1I/l
vr9Sn6QFZcehz445H5JCQ6SoDlq/NlJWBFqkDxrCnHIsQJ35ltng9307aD8veavK
oKYXM165+h8mxBpxSHIArvF1yd03BfJxMQI+ab82K4XrccyvzUdFzYK8srZjKpOV
MYNiBEJ9F8yCuMLfrhvja0VXxQpEVq+DYDGOIt6OuxVuKE1cMSPtq3IZLjimKpqk
/a9UNPjaybg7PFZzi8ArpEcyalUuNN+69Mcb10NBqBT3hp+a+ctSHqbvse5ff2f/
hFNYGJJWFejMRMz2D4TLx1EFVTQ0XmYwMzvskMXyYNQ54VvfosiJYLyYtiOem9kK
K0cgHaZ20YhHj6MeK1BwNj/mKtsmc9pDJb0gPMP/Jn2G/pJrIy2EaCNfCiBt+dHo
7TT3sKoICp7z6iuVNMgsgiGbLh4yUUecjA5/Ek+Ep23gJkxMcwAalxhBx0h1uWCZ
Al7qyWpKz5MmxjRCC5L3vtTHBgbC6tZhzpuX/vevLi1ezCFNHVfz8gwe9EK3GJAt
jHjIJsZQxXaLFaMselMlUMvvb5Yixep6Yf2F7NdVWBg4Qy4lVf5IQIwVysNLIQJn
pl0FrJVV8WS6/1BxMrDj/xT63xW6IB3MKL3IKDby/31L7bpBUWXdYlGJGxKl9bBW
gv8NY8Ru8vRyfTwPYffYWRnO1Iu54wkUksIBrOY6iiLJqSaBAP+fL4TMPlV8ZDPB
KuJJHUUmVM87TmEMsltP5PA1Tdixl+qdDDQqs5aC04SH8b3eMx0rFx0Xdf0UY9q+
v29PswW0XGKDvxN6SwOnbmYm21wLttBsD7Jig2kPmv4Jmt4uCVtsuvCX6wknqqy8
UyP0M393EQPH3T6CjzCQPUpOu4j4TgrS3/cQF5N2vj4lvGPWDBKga+EZB6msNKs+
2gny/HghcLIdmnwgoXNy7+dej4C5CnRzAoWCI3c9D7qqN4kQRPk/0itu9S88csY6
Wc7h5e9pdh2jq0pv5+/R5en3P29jvAMxe2tpeuP2uGBhtGL7WO8hL+IA3fM8sJpW
OVMhBP7tF/9RXuDVMIQRpRQC+CpL3JdXjqNl7qbdXiVxe6t+ESygTuXHLTbiX7V+
n+WxZeSp3Pk+tF/YZjanb7K3LN1qlPOsFl166vnuEVxf3m1Zjju78xq/unc3M4HA
DP7rAFuZcNfNPNZ1n1ygHZW4BKGyGeBEZMmptUfCIrSdmkzq3cZPfN2f3UHX2v3V
XqMw0KssWLk2lXe7NOCHLwZEAwTpz56640AkyW+kQHsgrxu0W7+Da+JaY4EWJpSD
0KC+kKOIE4SE06ucdw7DfccedYbvyh0fVbuUozzc8fXDQOTC3ZzOwsieep4idqPr
989Nm+PsGpoFkvG7bM/iq0yqZHnnko7DJqW+spcWM6nv1Eo8iX6dcTmmL8R/gCH9
m7D2uuI2PbpfzPxNe1h+8RmAzt9f0FOYfrQJLBq/DRzqHS1C2YOq+Lf/u+7U/PgG
gZY2fapZRHLqt25FWZxDSsZXVWdZf1Yl/Gv2lv3Q41U+Vy2hXc0+bwns3lvZMaPx
Rs1lHe1rafJBqLuP5RvPLgr6nipX2g0C4ONFDYHOF2GWOh9I6OY11XxzgM4kNqOQ
5hWL2YAhVXm3rvNu6CQGsUv56dwizvCEkVvD1Xt/Ffy6/2ZloTLMwrapOLhY60Dz
e5vCnSBT9LykQ0LpYYOxciVEkU+X/Ou+b1d5HFubZM5iJr4FklU8tLK4v8mn8IOd
qW1GIadJw8Lp8f+RNDrDPX6ejjBTgQqCC46GWdZtZS/4AVTGrb7rITDLB1/qR1SZ
23sDxEUbfNaR11SBzZXdta0A8dxj4J7DRMHSryGdU29bkirIIllyrvyKXOwEL5l3
wKseVXtBOFLWQxgF4NRzquA8zR/Hgarihq11obw9Mk2s8s9gqPsDuUlZJ8CIfp/0
WmwThjiPlxdHZw3VyeI4c+Q8sc7p+Iya2x7AKvpJfxHL2ecnaXgJQb9Ois3OCtiz
/q90xmeDSCFa06EPO806UbESlfDI5AE/lGl7nuCgYt/EbrQ0USEYe6C53z7bMu5/
PUvR218rELmVL42k/a6slNCYE7wiVsvABj3W72jhMHtE5o8XK335W3yZKqOM9NxR
GRME/f+PVPVdv8ykCUk5pLduBhxFeSoz1fzSwm/MC3lwRGwkxjvx5+ahPC+oyTMX
9lZqa/SWNmBgpPW7r4Wgk3Nw/QTAOdYI6BBo6tVx+IQ26yVAnFVmusXAAqPtspEk
XeLRs3ma1KYN3Aa3rCTIg+jLWPftSEjADPLa+1+AXDZn9XxXd1SEt9aKj+4Cfg7y
wkOV3kWfIHvrWozjZJbGmBX9PGStzzRzlQe0Dw91yx6GQ41GSfaXgmm9jrMh1MqO
5zmHs9SANP6SctFPB1gj0nyQJx0DiQ/0685C0eVVMDBHGZR6AR98xmDleXyBzkN6
YD9Tt0hE+dMLsImKU5mA/oaRFwZJJNV5lyfO4ofjkL9bd36rxt/iPbS4b/9FVdRv
dceQucl6ItwwsYSTjErE4HyiAPqR6Jp5azjpbTEmvTsRCsdBg2Da1Z2WmO4gtqj6
79MHngs3qx5O1QBa3A7thTJKjPObiaykAAzTUHTj/Lz+YGB/8B7ShYldG8o9AaKm
tEUjm7K4Ijaum5SmzWsjw8UrgJjsLzJN9rPdq1zQU4BPRlz79+pvXJCAfIEmXZ9W
a9ELsoB8POMrDIhsmkm6k+NcJc+zrDWUofKNG1/8l3qnaDDkyI5MRGOsSAe+bLWA
SlqMx6JzgL9noyjkG4vIk5Rv/oIvSXN0Iv00ejRZR2FuT9Ow3PsQsx3c2CVk4LXc
STfEx0Y83YR+nVFMxOojCm5VSnglfDLsA3JTWCrGd04bWv5TfQg1XJ0E9idoN6nF
CiliimXOMjTa0m9BtqwggifnzwOvWpPf16z5gZhHlW8/XIlcB3o1H2iH/1wGCxU7
Q910J6G8PR4gGaf6vQre0FCJsr5oR2/ST89xCFZ49ZUG4w9oBNWis8mUgmmrI/ff
iGcNChzBaA7pVSjSTD4sPssM+lLsgqAs/B8FQJbAUuq4xX96C3EY+X2fNa8KxF85
UdYeabOGYiKn5jx9AY3jLfpX142bfzy7aPt9nCGhJB9faLHNRZJHpQ1X8UA4QaR1
r1fjqGlCLoqqD7lTpk3fRZnPf7KwHhhL/BgvoaMbK6pmOGqsrIJrQHmP+ck6kUDU
2RmCsTZ3iRymPAOXGwWed4eCUor+xFR55ar1IohROSV+QRD2gzRof4Rrf0UJu2JA
OwHTC+fxqfWolma/kqyjN4wvD0Jcx6Sr1aVx+NDsZ18EoeOW23AAWssDWh6ZuPeK
uIwBFAwzUPl42WreniOC98mns8scUqVJPO5QfG97cet29VKYOxs5Vu4KwyPgGEtH
pPAhI981zBM7mmiVcIgQ3JC5lVmWXnqLjI9bVFQ4LlSi+LiDeoljnXh0gxzo5Ik/
Cl0Ho5oeDYCVCpPGVstfafr2Jp722dTxf90QTl7mArLW3a3MIX3F24bVvXAFZIl5
6nPtJP0mNU5lNGPwNe1oDWN7iUm3FBUnIDARhWUlNQX3UNlorREjNb/jm4QNasPz
eU4pWurMTjyOkCf9v7dyLeH/rw8ciSI30ojFTiJyP6E8dGfa2uVxngw2sQm1t2oJ
+TghHzzB8c+sCBOS5QXPhB9DRfktgOODUeGHuVb63NrzC374Nl+6M5xWuh/uS8Yp
GFrFoouVMLXRCi0tk1JSJSVb5ByV4iVFWgNseod+aSHbWc2eD0iGlTzgZd5Hzl+D
BH+4ATkvo0C8VGAW47RpTVWeNOmRB1KBD7inWVFL3+BtWXrejTz7Xk55rq5Vyddv
seSphjYoruLNW8lIUm/DEY5CWBzNZJfSsUo+VZWzMg3Vqm43xOmxOB84kTgXCuJZ
wEEgkYESoC6nnwALqgeIzlxBqkbKwTiIbmh69zFID8YtlchIluRqmyWGJi28IxNp
BdJxOHwOLMaQ2SXBevBqWk9nhZczmg/IBhVbihSk1Yu+4Wlp0ZAB72PhaElbBnxt
kcz2NLsVV0Q3ZPh5kJeCWLsOFR65j9eKCyeSRn8rUHxuSM+jlzOFJ4dOS4+WNG7E
H4xKFeFCW42OX78t2GSX1PhwCKWhGR2CUzAlYkvNDgJP8jjLy6PxBri74NGIWo9L
jRqJ5/IQOUJBOVD3iYUej9Wz1K8QGfxxu5FtdlGI+G+DPuFp4UO2D2p3znnSz+Qt
bU1+vrflBAm3FBojritn+sJwa6yeSfiGOy6gCQZX45LiL+42+AUYJFudq+ViW6+W
adXdSivJI1ORURzp8RQLO+geYT45THAGsy6LVjvOl7FHttvGgNZ9PLAnVc7lZc33
dpCsBP2X/LaQnjRM8jzBm5YWCXN4V5AdCY2qpzqjpLxUJHGhmHY5I8xerA/VvgjP
k9vguRrcyzhtt6igX0+9XZwFZKNvJxqq3ewgmM6dwIp7UqGwjFCV8mSKDYS2ciP0
jO9Mf//YEr7Wxr5UzZo14r9h2O/2b4xgQKDTiPmZX7u/abJ4tR06sJ0EcGeZLVSc
GKE6BEheZxhHAovlfZrgZRPFiImYemj+OLKx/54vE8omlq0YgbS6m9xf6qUqQZo7
DOvxjCnmw6pBv/gPOu4z7zSK0I2CIRYUZxZsIl8sWNif4/sQeOT97bgkN+lI3Ln2
obkGtlVdGFnv1sOLcxXLhU9qtiDXt8jlCm8IMA3fFs5qzLMhmsRNrf45Z/eybXSX
XPCK0LlN3uRP5sttwwBFgiLmznBLsSmvwFpYDe8NiALwLRPLthyIUXH71Nvf1CSg
lae3VTOvuyyDtIkoAaOz9UV9MlLwmfWDNBgVw8OpcUo/uRU13sF33YRPXLyDx1Tc
sQX1Pd9rptTe7KpPZ1DijEvpkBZupvgJ7zwQyZ5wUu99GJTI1bjyahFdAtEFUNZZ
/FeXJutxAXV3oIezRyblsaZO4xNizvLyDANZL07wjHk3jBM8uy5xsI3Gcm2x+R7B
p31Nb8pq+667Bm8B6KDxzBsToJaxMrM03T3XpRaDt+CZnVERAC6I686ZR6oYzmuw
N5lCjxr6W2SUHK276/k3cX8Nuudu53p0mrrR87ur5IwgwE/AwKyoLiYMZHZUcsMy
zn/4vC0MCSEmjcCa4LFVUOzEsilMHS6eEn/mfKB/cD4gfIggjH4QQHaO8ipls1rY
IyF5JbS9GLzvNOiWUhmBHPVP9R+XCMZOBi9lLgUUuXf21/pJjnkIpH0LEYLwkO4A
qL3Ci8UPesK4eJ0vhjDhf4bhlrZ8hlUl8dDq/n79ku9ctBDbfo3zqfPPRoR7g0O9
jNkuQE96YcoInwOBflZ/tUaN1+u1v2VA/wVKQng0CmWLRaRg/+0sUCbNuzxSJEBk
IEofWKNKoxM7fBoaeMnz1JgayB1gsTA3EUMZ7DL/Hhtm404HAXZEb2rr5xHBEMaQ
fYXCHm2mbjxm0QIy4Uqc/MFUzRd+RgWZ/GxdGBRFLjnedwzMwEAiM3sy0BNq9lAh
9fEIcnYPQXQuJ+qpr1DeWTbJz9vGlyzWl0FW3QBgWeyYn4BrbGQzMy9f9t86W4cf
gWBezjEbbVe5V4sTJH76RSkK2qIE+0DqMvW1Qm8ezBhQtb9YVbRzOn5A4TKuFdLv
jltwSHH1xJlPieH2bak2Cm3R7O0MFq9ODpKh0xhm7PzDClUKa/JXmePD0ule23Zf
VK0jgvaKTIsgQAvxzFdLm4N4G/ZJvIswKmYlCiKw9N5yMUZrXWCSrcnM/eFDh2XA
zabIohdvCsHfPoeLIJj6gwiTNJ26v2MqvximrBDfRuaGoEfUkbAWbwysKGOPbeyX
OGq4foBD7w9XxXCmwJ0BLOJKuRwl1GKTYaaqLKC8Mc2CKllgmtRIJ1n/Q/hZlXUA
7+qmgpf0e78KZxnLIVVG5UnfOet+FcNVeB1HKUZDHtPmy3sHs1JL/moJ0iWNYqbv
7OCCSgWgZ9+161z3E0tGQSOZASlQ2nHkfhOa68BaKx2W3GG1h08cQyiquc47C1d9
plEaEJvpqjaQT92XHMHTHeqLiDCU68wz4pZ+EOOQjUZBRDa9QYINfQVI0JMkWGUF
ngZZkK0qeaJxridBA9M/zQqKhW3Bmtm/90nRKbLyEDuqdfRdXfgkcpFbE7b39Ysf
nAgVfO37gMwRtNFaAfQawyWH9hetkjV2u/KQt2CHainpKpbdiWtBl1NFTtZGK+bl
eQ3P4nCnKWRZNK+GKSOYndvNxMTyUGg5NGUv1jTvwY4SR7b5/Ei5YLjlHTJnOw2d
8uvxTGmAb/5jsV0onYMkLQfKxOUcypu4bJFojwdDE36Qb+ZJtu/59reIHFnulGrT
4ePegYuGpkKeu8fojvzbzRsI6889nv3rtilQUQW+NqQf0SYXu1PoUFJ0GUJBZh2B
9wWgKFucVdekQPlwzvKInxF7v5KU0jTwfWAcISn0gKy4IEzIuWPltPa14lEzoIfu
m+VWej/qGbKW9GyfhShxkHFO72ci9vulDn6T6mriNJ1pLChtkg9PVnY4bY72d+gm
NCFzKwLbRERdK86weFB5jbwny2bOWJcigRbr61h8R71TvGABCVnTCNS2ssGCPqRQ
8nha4xNYixpF3jB4gQ3hFo6Ukl1qkAkyhtYJptlshUTLimIt5JCnDRNEb6GhMGq7
UKi6mpTlamumJ+0hMeJBlWK8xRce+Iy8LriJDqfz07bqvHQ580ZAce5PyYNlOEDS
rCTremE39Mx5Cy8iMNJ2UQtTEVKX82RPyca35zpD+HAF4vp8vpZpg7+owoYz1wyU
Edtry8Ojj1s2DpXa1d+FChhA43+5wylj/OmAoCxhMoxVOBNobMszpYRQ1vUrmioR
PkmHMnScclmwn8iUHaDiTAkoQbB8JDeiZFhJPGUJpURgQPUB8J8MILEv+9X9Pb6F
NUklJ4Qk0XknWnrJUE9dS7fiUp6pATLGtgTPSg2McBjOcotVZugED/WjPWSAyS+6
O8cCl4TNigidt/S3xxv++w2Wn4axYcM2lDqmzSbK+axZADY6Lfl2aFc+XGbI5byu
oJNTvNHn2NL4BT3WHZdLm4MhheTD+9JKOI8afd1xAxs7LjXWqYv8/jM/UGXfECLL
IE3Y6w/+TWOqRypiVo3owHwq7RtMpVS+4KrXEva1EIZT3CLsTU+Njf3amtapeN4Z
PR6lZNCZHIXJTH+XrOq+6N+t/IKmyCM6fk7xFtX5JMybRdOk07HSIjiOw62/BiPv
Wr5xzPoUI5z0VrM63Rq3EvhxwXAlNbCuTk64nQecGwJWG+ETk9no/1rdi23NkhfB
+p1N5bqquFGiSgg4EdfeFDVqQAI2HTIaqId8Mw8okQbv6N4u8jTf4+zv2TMzM1MF
TwbPiKJz3lTbzURwnQNJl4etE9iBG99q29/DFamo5VD3JUVLTCmg87H9wc/xvCQQ
4NfmdOBO9ypCZ7odHpBPKCwni0xLghFcyIhbpv/44imepi5ZL3cENBELwE0ZxDJv
3Me2I0+btxv0GajOjpvaEutUFtaNpMyi0AobqEWhVuTCRNIYQw/IosPT+DZDQVaG
zm4B/Xwqf1KdaBytOJj82UVXB5BFsy22PL3aa+H6NVnWUN5Z7pTrYFyiYjoJTk+T
d7rJ9kUqluZ+IsmU2/+xxFgBUu7qTC8wEThWAzJimQ11tZmSZxb8dTyeeWHBL5dI
4ycSiq6zGjUUdofdF1BoQ5mt+Q/cUl20kljTYlS2yZnkk4jYd9tK0WbSn1sl1QnP
T7zBYwUSgaTsUV5ilzrZ3CSDr8i9ykd6Rj+Chs9B8S03FSoBCBUJr5mYjpSw8X55
hCDBc1NsHZvXu5Yg08CrsSuqGCHCv+fnJU0P3bthdjUJRV+8Zb9XnHXsj/LZDqxG
XguilICEgSjGT/ABmlU8PfCARGbNkl8wsESoGQJm7JQkTLFHlN/cC5cGePjk5i7W
c/xod0SmRA0qrwnC6ZIXoyOdn91OFsikE2PpDJN/aBNC6j05p2RgwEzd5gy00ueS
WH1OwT/ve8blxU9P6Sq6/DuIdirgCpIDW3eTyTgm6Yt4R/mMXjDURTiQHW6f6Ye9
6PNvKuBBVGDMiNUmWc3gB/mvJ43UjcDOGj74S9A1sYUflIy1jmCz18Qb6yskaNBQ
CNSmka5t4hC/5JYTfuiR0lWiTTcRwhJMi3IKp3kw/plvvRQ3jsXNsQbAOBUfEKtR
Zv5wT2B/kQRnXT/NYJnnpv0akR49379zNldgexFyHaX2ESpV+m7Efdlmn98mNJ5u
DJm4v1FPDULSbNhPHTPc4NdxHjo/IY4WNVz6JiG59h3L0UbJzLOCziwSTsoLihIU
NxNms/2mAOKtCwsUkTz6jOUA2WLLAlQ/fF17EtmsrI2UtcqE4DFYwMH4LxDIsitq
2n6WcJ1QTUHdynDPIeW9hI3Jcx39k0lNKIcDx7c2DbXKqLFsBQY8mbrHJfJ7MduZ
KgnCh27ZhLeCht/du/lfA+yZaRhycr8llDpZVztnB2tyUqMEaGgu5GJSgJV6FmFK
VfKHNlt+8wP6wT8GqJmdtMODdm6m3/oAX3Tba3UxU5gyHu+kQUNTNOiC89Nysvwx
wkWoKUPkEYNBf1o7UT0Ywkc1ljmxXfbLXHd2Lsn8ZEjy6A9lhNot+qvze/d0IV/b
EVapStrKtv68hq8Vxemrdvszan2plP9v15VuF3mBEqisgzpptGL8jnKvUP6QHvG4
rJt+4JWEHC1BN7dOETcEDx6vt2pYncmKs7kRBvWMORdn4DUJrrwIcDx20wc3wG63
+VCCUZtctcl6oGC+4SUAdGNEan7JeVif7We//BAyZbtvdkkL+Kge2rsW9Uq7vJFB
8Rbc73UMseuZI/QXLtOjBhS4PrmPTG1F4f0kCRb5ANaoUi1JiQVvhqOLuTmBk63t
32Pc9S+3QHJXK/m5ryy2MQ/SyoDlDkx8leaNKJ231LFJXkoqqUdCDyvwTTf4dWx+
FDz2dPawHcc4Fc39AgBHKA==
//pragma protect end_data_block
//pragma protect digest_block
SFGH+WKKoB0m5pX7GREaHK+Wf2I=
//pragma protect end_digest_block
//pragma protect end_protected
