//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
84MC8KkO/kry6BqVXmzUHmtQzlB2JkBnMDunX0NfIXqaTBdaBBVdK5vagM+cbGTs
Qu0LYiaRcplI9GVzJdE2P7ahJtVxEzgT6TAbF6Bl8bBunHbROx9oSr9HnGsMwUZe
1wElfMgGEWFRnKA2XVbebOybWQMo/MPZBq1pP9QH5vu1nXiW3tVmsQ==
//pragma protect end_key_block
//pragma protect digest_block
dCrsjeyV7teoJjWChrDln9b3RB0=
//pragma protect end_digest_block
//pragma protect data_block
Us4wVTNyd7NEMOh5ngR0YCrk0hF/FwrtHONBvCjgY6PD2bHBVFG738OiGUJJ3+gV
mG1NRD9FzK5619aRpKpsBkDqO7g8W1EL9INzXydiLBwOTBtQyqNglmYe++l2jpgn
kV6teMQPgnWr3T7sdY1+Va/BZlvGCcOoQ7xwhkPHAoaC/x8o6Dg690XAmHw+Q6cC
yTDNgJOL9XeUeu26U+3CzmYw3+d+F+E44ZdocAajtDe7UJhBZpMSMzfZ9vmFd4Iq
D73fIy6Mq0PHWA0CL0PwMDqGHOE93vUPWmJWkwBfQ+t42UQQjSQBLyH58JmvZ86O
QxCblNR5Z91R2Y/qSiPXzE/HhthIEHxRhtYvvDfjUtfmAg/8/Uy5lQUtrAPbrvqq
WgQQKlwiYarGNNXRh+qbwRrHT8asMTn/YOD/iA9VLqcvIWdE0gTDVNImZkhN93s1
RLBl2r4wynozQCO/QQEma2d0/IK/barmMhVvqxg/J0SnRfyiuu0nA8+hAwayZXGe
3EJE32u0hJ4/801vT1Iox/n+Abgu4mmF77C3+gMmOaSfxczI0e5YsX6Zj2L47q9a
bO5OFls6E6/eoqTpDnm7WLpop1NigwfXih9yD01bUyfIkntS0b/rMB45ILxSScoC
LSlNukK+bGALwKEx9hvWx+ZQuG8jsGF5FXXgyVmB/Swofsb0B+nytvWjNw++T96a
vhxUUjupQQIpjT0+aUXS5I2ygN4u91WiYX2Q3M0OovXKqeN37dUysK2Vh7lfKoCE
M3mT848dUof/hIPBqh5pGEn5CiG0+qqr1pqjNsTK7rQh3rJbP5wFm1XMzlA6FlMY
LvwFa+XEWr6rde5W4H+QRP0Sv34QNDvFptCgG/NntCmHQc4siStMlAs98mwTQeMJ
tfLZZQy7JqQ4dlSV9n3LyqmdMOLQCopbol4RrNBtTaQfz8Yd22eZ0l88oytA9lcC
SQL1lZ7rdi9swKfIXZ+cgxKPI9smDPvG7bfupNSwX53FwQ90DC4lyBK5Lv4N6p8h
hj2wemFF/8iAI9uSebZF9iCaCoHPiJgR/sYi/zswpVFlpOp4vXWd5upSFe379q+o
WkAduOFmjNeHuX9Cuqi2DtQ8uOWlttoV4+QoQpCA337R4Eet+KH5mVUtdqKlMv8O
1OcZsssOQ/9e1t+QpHyWgy4GUZgJfhOkASeuvbGf5+C17ZvynfNJMJHIOI9fAnoa
liyRq6pc34RanEOjJYmj06lj+8yE2E7Rwzi8MfgxrbjsQZ9Gcuafq32O+7W9PsZx
3KQx/bLCbwtyqOZPz5HA0WY2litzHzZhchaUZuqya2NOVShuXw3NvZTC+ykY39K5
2YWib/8A1rlD3uoy3oMRePao2GB52zNZkti60n3k66uDknX2Ft9hYEr24Anxv9P2
JIgmk2C5PxRt9QaCnbspYKJeZxL7DTXEtRzgJx+rPhk2e3bE+YPY3aCGpziErkg7
+nOszX6ubJhj+eQ8TlNwiqLKcX0tZXcuGCythCOg/9zVqOS5CvdJa1Ki02XyiJP/
Ibua1cNfXyJRapM83/SCv3IPSziGjm+6oo0OWMQDiJaCMHxq6VsomRXlWuLsVNY5
4dZLwFmJzOjMw+4UDyv50ip9l3Mm5N/3U7mEpDh0pT8a09DwrZBr0yrkEchr4yzg
wvbvHiveDheGCX1pdu5JwuzsmFRiz/d23KUXUweR2soUZs3FCa/widAluMX7Hvw5
nckKKsKzlPH8RTpsLPy1IjOS1gpYfJi3Kk5Q10hY6FJE7OQi9jOaGP+FYZ2XzZV6
RB6Y2loPdAM66jL0JrLzWZ7qWUlNJfHFULtLy6als2EXnk/rk9KbR0gUlpnSUolo
oRkvE7LMQ2ICPniVkX+lYW4+yMyhDKf8uBKvVOXYl2pvzwgWrhFuUTlvh4z+ygAl
XtQYTRsZPNpF7I9hz9CdwL1H50yBam3UM+eabrqZsk3uyDD+VvbzHQfZivGrfiqJ
nS0SIHSefAp8aTnSsi7NnPAJlwA/QG9g1us8CFe6vv1U5/wDOqjrWYpJ3AaQSdfx
DwLJ1JzznY76UMgSMv+HJTr9jgSpr3llpJz68raJNurOacDxXqPaYOyd3a65JHpE
AxVGDkvrt0Sc0TB02FoaskbgR/EofSRR0qQOymYGHR5RbjlAQs5yjw0Ljk07LiUx
sYSjmJ2wDwCXQ6MkukLvk+K2MoPELcQU06YnnDXJOfc/qHAV8pipnZ6PMkDq206P
htzYLgo+yYiEAzQHDyxhjMTNRTbPl62PZnIVqtJa1WXq6o+PKUcWFtMFnMpUDNBr
aNDTuhukC1ieJnHp0MAzKjFZEmg79C73k1j7Nc9RpyNqKXzs6jhwl9On99RIAknv
Z4RqtpwXnANm3P1gLdsngZSaOiBUTqBLqOsyQcmHyuxUSCg1Yoj5RM93qvk+leBo
rXApLggNmvl/+0hwaKxRqpZ/7AJQBNcA+F9g8EHTG1tbWg6Lw5P9GJSF9SCAvIZv
SQ1sEVQiUmPgSpG7PlGt1LgOMwVSlLs1sMJ8Sthu/5dK4PlVoeTQ1SNbtsEmVSQp
/AIrwOrAsbVFvruRdM2s9cD7TZ5wYQ7uRZ4loZkqqgN/N3jWxmq27+nBQvKdiHZe
wplTD/YTIuPXQ/PhbMHnr0mytO1AUwVJ13OzZ1VkZqcRRbeR9ZHlCHIan78VnEwQ
owKn7QBCu6zrXaRSDSYPDI1f8RJSUEBvsJMHMVOMgSA6/kAoVfwpdZMnK2nw6WbS
Ir6ewTKMCprQZrGth5jAQU5K1ewBclh/GkO91xw5MEgTfZAa+oSfI8/Z3irgY6e2
bgGypmvKWfR4z7O6ey6bh4U5aegDygWkFTF92RWqPOw7X0QLLNmffXS+dNA5ZRpO
F3ngTILVLDUcn92xeTzXhtCHl3Vr2YT0Yl7JC/S/jvu+dHNz8dpo8Y1+AhNn1/le
iJ2TwbyPx3YNGGklmzmviF3KWEF+21M/T4TvRWHJdb3oAz0bRbpDaRLWkNTiGe3I
5RN6vjt/gX+MyMowPFpjte2UqLcF1sStLeSozd2KhYkuLOGRoeLLpkooI2LMvjIP
qkO/6CYAK5uoe3MifhoUOh9EVFugZ+e6K3M0ELAQhm3bNg7+C1dSFbk25U9lsPHD
d73qaj9pvmldbXk9eFI5KBfD543mJjXeyBuEzW4yi4VPtEV7A/WyFPOpnZIoMGxw
KXsNvFx9QvWwi4NKnkE17MMIuw00iWvgFVFjK0Rik/2slFHq3k717Xn8XcxuKE9O
3SvVrufp8MbE8hVgiDVc/DJeYlJ4n4KIPiFV9AKZQF7V9n7iSRrud/wXL3rmFIWa
gxL/Ecgj2gpWd6mYw3YrlsRsNZDVULqgKJrfKPctaiotelP0iV/5oml1OWxT5rY8
EFIs3fx4EFH0ADC4wBZMEMN+bDWuXSzPXa/wr0SAruTuQJYKuEdCw52ikbVzt+6I
NNreWhsQ7TDyX0AAsq8BF/ujE8+WOy+kCV8kns/HQLi7HOEfGUpimSQHa4cfHXQp
AlMe0Y7isf0tiI6AyiooKeC3bE9DP1SwQaGT8TcNksK1CWC1Zf5f7551ovzHgfkl
rfXAdpu3oPP6xjY7Pkxkfq5TMmaKlS0U0auzyVnLHl0SbWMLqMeW60Ur6ECiBHR0
07+EAAp/HuvqZr1DFBv6LyMEalo8YrhsgOEIJrlyB9081+BDMKhvIZxD8oF1Adlb
9Mo/ihiozR9KRnkQAZhLZ1t5WsoQ+n/eUoRCGdKcjXfoF5tpKXANKANe+JSJ++NW
YqS55WL4WMkrDpgBs6HP+2xCioNMrEW1/r9fE+fFQ1tXBylD/VN1ePbPD42tkcHj
DY235mc3ktQez1FzG+yF/0bti45XG9dzfWNIrcVHIz6mqe30QEUKZRPh98TCCH42
5NAYPmpNo9iVKqMUk8LFOY2Sg2aS8E7cjUnFkqZrzjV9zlmeMWTQdymNffYKUy6t
DHQFTUEKUprwgCSAi5El24P/qUZ8UA6N9BUCZyjKf6wm8tMB1Z1031mSu48cUb5k
g/7mWHciVEqeAtvAueAfR+agi/V4b1qFO4hItiIXWke8EaOJpiVM2ZAiaoJ/Mrem
juAF8Nx7UTs7rZi8xhm5HiPj2sfcX0EDBt3eNGof9b5skbAzvlqoFcjvoFl2/X3B
yWy/LQn0MX8+RJMbkTrWDnsPS3Thhpb1AdvhKaRVvLLrgiePvf8eFTD2eMVqK2Bj
577+IGbFd6Iz0EUJ73b+pz1bd34oLyaj5WiqQKEYOKdTOy0jtygqlYSXvqaqm/B+

//pragma protect end_data_block
//pragma protect digest_block
Zmpkfa5WU0/YHbuYVuYtvoJJFfQ=
//pragma protect end_digest_block
//pragma protect end_protected
